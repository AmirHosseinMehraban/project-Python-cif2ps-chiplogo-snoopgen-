magic
tech  scmos
timestamp 777777777
<< poly >>
rect 3 64 4 65
rect 4 64 5 65
rect 5 64 6 65
rect 6 64 7 65
rect 7 64 8 65
rect 8 64 9 65
rect 9 64 10 65
rect 10 64 11 65
rect 11 64 12 65
rect 12 64 13 65
rect 13 64 14 65
rect 14 64 15 65
rect 15 64 16 65
rect 16 64 17 65
rect 17 64 18 65
rect 18 64 19 65
rect 19 64 20 65
rect 20 64 21 65
rect 21 64 22 65
rect 22 64 23 65
rect 23 64 24 65
rect 24 64 25 65
rect 25 64 26 65
rect 26 64 27 65
rect 27 64 28 65
rect 28 64 29 65
rect 29 64 30 65
rect 30 64 31 65
rect 31 64 32 65
rect 32 64 33 65
rect 33 64 34 65
rect 34 64 35 65
rect 35 64 36 65
rect 36 64 37 65
rect 37 64 38 65
rect 38 64 39 65
rect 39 64 40 65
rect 40 64 41 65
rect 41 64 42 65
rect 42 64 43 65
rect 43 64 44 65
rect 44 64 45 65
rect 45 64 46 65
rect 46 64 47 65
rect 47 64 48 65
rect 48 64 49 65
rect 49 64 50 65
rect 50 64 51 65
rect 51 64 52 65
rect 52 64 53 65
rect 53 64 54 65
rect 54 64 55 65
rect 55 64 56 65
rect 56 64 57 65
rect 57 64 58 65
rect 58 64 59 65
rect 59 64 60 65
rect 60 64 61 65
rect 61 64 62 65
rect 62 64 63 65
rect 63 64 64 65
rect 64 64 65 65
rect 65 64 66 65
rect 66 64 67 65
rect 67 64 68 65
rect 68 64 69 65
rect 69 64 70 65
rect 70 64 71 65
rect 71 64 72 65
rect 72 64 73 65
rect 73 64 74 65
rect 74 64 75 65
rect 75 64 76 65
rect 76 64 77 65
rect 77 64 78 65
rect 78 64 79 65
rect 79 64 80 65
rect 80 64 81 65
rect 81 64 82 65
rect 82 64 83 65
rect 83 64 84 65
rect 84 64 85 65
rect 85 64 86 65
rect 86 64 87 65
rect 87 64 88 65
rect 88 64 89 65
rect 89 64 90 65
rect 90 64 91 65
rect 91 64 92 65
rect 92 64 93 65
rect 93 64 94 65
rect 94 64 95 65
rect 95 64 96 65
rect 96 64 97 65
rect 97 64 98 65
rect 98 64 99 65
rect 99 64 100 65
rect 100 64 101 65
rect 101 64 102 65
rect 102 64 103 65
rect 103 64 104 65
rect 104 64 105 65
rect 105 64 106 65
rect 106 64 107 65
rect 107 64 108 65
rect 108 64 109 65
rect 109 64 110 65
rect 110 64 111 65
rect 111 64 112 65
rect 112 64 113 65
rect 113 64 114 65
rect 114 64 115 65
rect 115 64 116 65
rect 116 64 117 65
rect 117 64 118 65
rect 118 64 119 65
rect 119 64 120 65
rect 120 64 121 65
rect 121 64 122 65
rect 122 64 123 65
rect 123 64 124 65
rect 124 64 125 65
rect 125 64 126 65
rect 126 64 127 65
rect 127 64 128 65
rect 128 64 129 65
rect 129 64 130 65
rect 130 64 131 65
rect 131 64 132 65
rect 132 64 133 65
rect 133 64 134 65
rect 134 64 135 65
rect 135 64 136 65
rect 136 64 137 65
rect 137 64 138 65
rect 138 64 139 65
rect 139 64 140 65
rect 140 64 141 65
rect 141 64 142 65
rect 142 64 143 65
rect 143 64 144 65
rect 144 64 145 65
rect 145 64 146 65
rect 146 64 147 65
rect 147 64 148 65
rect 148 64 149 65
rect 149 64 150 65
rect 150 64 151 65
rect 151 64 152 65
rect 152 64 153 65
rect 153 64 154 65
rect 154 64 155 65
rect 155 64 156 65
rect 156 64 157 65
rect 157 64 158 65
rect 158 64 159 65
rect 159 64 160 65
rect 160 64 161 65
rect 161 64 162 65
rect 162 64 163 65
rect 163 64 164 65
rect 164 64 165 65
rect 165 64 166 65
rect 166 64 167 65
rect 167 64 168 65
rect 168 64 169 65
rect 169 64 170 65
rect 170 64 171 65
rect 171 64 172 65
rect 172 64 173 65
rect 173 64 174 65
rect 174 64 175 65
rect 175 64 176 65
rect 176 64 177 65
rect 177 64 178 65
rect 178 64 179 65
rect 179 64 180 65
rect 180 64 181 65
rect 181 64 182 65
rect 182 64 183 65
rect 183 64 184 65
rect 184 64 185 65
rect 185 64 186 65
rect 186 64 187 65
rect 187 64 188 65
rect 188 64 189 65
rect 189 64 190 65
rect 190 64 191 65
rect 191 64 192 65
rect 192 64 193 65
rect 193 64 194 65
rect 194 64 195 65
rect 195 64 196 65
rect 196 64 197 65
rect 197 64 198 65
rect 198 64 199 65
rect 199 64 200 65
rect 200 64 201 65
rect 201 64 202 65
rect 202 64 203 65
rect 203 64 204 65
rect 204 64 205 65
rect 205 64 206 65
rect 206 64 207 65
rect 207 64 208 65
rect 208 64 209 65
rect 209 64 210 65
rect 210 64 211 65
rect 211 64 212 65
rect 212 64 213 65
rect 213 64 214 65
rect 214 64 215 65
rect 215 64 216 65
rect 216 64 217 65
rect 217 64 218 65
rect 218 64 219 65
rect 219 64 220 65
rect 220 64 221 65
rect 221 64 222 65
rect 222 64 223 65
rect 223 64 224 65
rect 224 64 225 65
rect 225 64 226 65
rect 226 64 227 65
rect 227 64 228 65
rect 228 64 229 65
rect 229 64 230 65
rect 230 64 231 65
rect 231 64 232 65
rect 232 64 233 65
rect 233 64 234 65
rect 234 64 235 65
rect 235 64 236 65
rect 236 64 237 65
rect 237 64 238 65
rect 238 64 239 65
rect 239 64 240 65
rect 240 64 241 65
rect 241 64 242 65
rect 242 64 243 65
rect 243 64 244 65
rect 244 64 245 65
rect 245 64 246 65
rect 246 64 247 65
rect 247 64 248 65
rect 248 64 249 65
rect 249 64 250 65
rect 250 64 251 65
rect 251 64 252 65
rect 252 64 253 65
rect 253 64 254 65
rect 254 64 255 65
rect 255 64 256 65
rect 256 64 257 65
rect 257 64 258 65
rect 258 64 259 65
rect 259 64 260 65
rect 260 64 261 65
rect 261 64 262 65
rect 262 64 263 65
rect 263 64 264 65
rect 264 64 265 65
rect 265 64 266 65
rect 266 64 267 65
rect 267 64 268 65
rect 268 64 269 65
rect 269 64 270 65
rect 270 64 271 65
rect 271 64 272 65
rect 272 64 273 65
rect 273 64 274 65
rect 274 64 275 65
rect 275 64 276 65
rect 276 64 277 65
rect 277 64 278 65
rect 278 64 279 65
rect 279 64 280 65
rect 280 64 281 65
rect 281 64 282 65
rect 282 64 283 65
rect 283 64 284 65
rect 284 64 285 65
rect 285 64 286 65
rect 286 64 287 65
rect 287 64 288 65
rect 288 64 289 65
rect 289 64 290 65
rect 290 64 291 65
rect 291 64 292 65
rect 3 63 4 64
rect 4 63 5 64
rect 5 63 6 64
rect 6 63 7 64
rect 7 63 8 64
rect 8 63 9 64
rect 9 63 10 64
rect 10 63 11 64
rect 11 63 12 64
rect 12 63 13 64
rect 13 63 14 64
rect 14 63 15 64
rect 15 63 16 64
rect 16 63 17 64
rect 17 63 18 64
rect 18 63 19 64
rect 19 63 20 64
rect 20 63 21 64
rect 21 63 22 64
rect 22 63 23 64
rect 23 63 24 64
rect 24 63 25 64
rect 25 63 26 64
rect 26 63 27 64
rect 27 63 28 64
rect 28 63 29 64
rect 29 63 30 64
rect 30 63 31 64
rect 31 63 32 64
rect 242 63 243 64
rect 243 63 244 64
rect 244 63 245 64
rect 245 63 246 64
rect 246 63 247 64
rect 247 63 248 64
rect 248 63 249 64
rect 249 63 250 64
rect 250 63 251 64
rect 251 63 252 64
rect 252 63 253 64
rect 253 63 254 64
rect 254 63 255 64
rect 255 63 256 64
rect 256 63 257 64
rect 257 63 258 64
rect 258 63 259 64
rect 259 63 260 64
rect 260 63 261 64
rect 261 63 262 64
rect 277 63 278 64
rect 278 63 279 64
rect 279 63 280 64
rect 280 63 281 64
rect 281 63 282 64
rect 282 63 283 64
rect 283 63 284 64
rect 284 63 285 64
rect 285 63 286 64
rect 286 63 287 64
rect 287 63 288 64
rect 288 63 289 64
rect 289 63 290 64
rect 290 63 291 64
rect 291 63 292 64
rect 6 62 7 63
rect 7 62 8 63
rect 8 62 9 63
rect 9 62 10 63
rect 10 62 11 63
rect 11 62 12 63
rect 12 62 13 63
rect 13 62 14 63
rect 14 62 15 63
rect 15 62 16 63
rect 16 62 17 63
rect 17 62 18 63
rect 18 62 19 63
rect 19 62 20 63
rect 20 62 21 63
rect 21 62 22 63
rect 22 62 23 63
rect 23 62 24 63
rect 24 62 25 63
rect 25 62 26 63
rect 26 62 27 63
rect 27 62 28 63
rect 28 62 29 63
rect 29 62 30 63
rect 30 62 31 63
rect 31 62 32 63
rect 32 62 33 63
rect 33 62 34 63
rect 34 62 35 63
rect 245 62 246 63
rect 246 62 247 63
rect 247 62 248 63
rect 248 62 249 63
rect 249 62 250 63
rect 250 62 251 63
rect 251 62 252 63
rect 252 62 253 63
rect 253 62 254 63
rect 254 62 255 63
rect 255 62 256 63
rect 256 62 257 63
rect 257 62 258 63
rect 281 62 282 63
rect 282 62 283 63
rect 283 62 284 63
rect 284 62 285 63
rect 285 62 286 63
rect 286 62 287 63
rect 287 62 288 63
rect 288 62 289 63
rect 289 62 290 63
rect 8 61 9 62
rect 9 61 10 62
rect 10 61 11 62
rect 11 61 12 62
rect 12 61 13 62
rect 13 61 14 62
rect 14 61 15 62
rect 15 61 16 62
rect 16 61 17 62
rect 26 61 27 62
rect 27 61 28 62
rect 28 61 29 62
rect 29 61 30 62
rect 30 61 31 62
rect 31 61 32 62
rect 32 61 33 62
rect 33 61 34 62
rect 34 61 35 62
rect 35 61 36 62
rect 247 61 248 62
rect 248 61 249 62
rect 249 61 250 62
rect 250 61 251 62
rect 251 61 252 62
rect 252 61 253 62
rect 253 61 254 62
rect 254 61 255 62
rect 255 61 256 62
rect 256 61 257 62
rect 282 61 283 62
rect 283 61 284 62
rect 284 61 285 62
rect 285 61 286 62
rect 286 61 287 62
rect 287 61 288 62
rect 8 60 9 61
rect 9 60 10 61
rect 10 60 11 61
rect 11 60 12 61
rect 12 60 13 61
rect 13 60 14 61
rect 14 60 15 61
rect 15 60 16 61
rect 28 60 29 61
rect 29 60 30 61
rect 30 60 31 61
rect 31 60 32 61
rect 32 60 33 61
rect 33 60 34 61
rect 34 60 35 61
rect 35 60 36 61
rect 36 60 37 61
rect 248 60 249 61
rect 249 60 250 61
rect 250 60 251 61
rect 251 60 252 61
rect 252 60 253 61
rect 253 60 254 61
rect 254 60 255 61
rect 255 60 256 61
rect 256 60 257 61
rect 283 60 284 61
rect 284 60 285 61
rect 285 60 286 61
rect 286 60 287 61
rect 287 60 288 61
rect 9 59 10 60
rect 10 59 11 60
rect 11 59 12 60
rect 12 59 13 60
rect 13 59 14 60
rect 14 59 15 60
rect 15 59 16 60
rect 30 59 31 60
rect 31 59 32 60
rect 32 59 33 60
rect 33 59 34 60
rect 34 59 35 60
rect 35 59 36 60
rect 36 59 37 60
rect 37 59 38 60
rect 248 59 249 60
rect 249 59 250 60
rect 250 59 251 60
rect 251 59 252 60
rect 252 59 253 60
rect 253 59 254 60
rect 254 59 255 60
rect 255 59 256 60
rect 256 59 257 60
rect 283 59 284 60
rect 284 59 285 60
rect 285 59 286 60
rect 286 59 287 60
rect 9 58 10 59
rect 10 58 11 59
rect 11 58 12 59
rect 12 58 13 59
rect 13 58 14 59
rect 14 58 15 59
rect 15 58 16 59
rect 31 58 32 59
rect 32 58 33 59
rect 33 58 34 59
rect 34 58 35 59
rect 35 58 36 59
rect 36 58 37 59
rect 37 58 38 59
rect 38 58 39 59
rect 248 58 249 59
rect 249 58 250 59
rect 250 58 251 59
rect 251 58 252 59
rect 252 58 253 59
rect 253 58 254 59
rect 254 58 255 59
rect 255 58 256 59
rect 256 58 257 59
rect 283 58 284 59
rect 284 58 285 59
rect 285 58 286 59
rect 9 57 10 58
rect 10 57 11 58
rect 11 57 12 58
rect 12 57 13 58
rect 13 57 14 58
rect 14 57 15 58
rect 15 57 16 58
rect 32 57 33 58
rect 33 57 34 58
rect 34 57 35 58
rect 35 57 36 58
rect 36 57 37 58
rect 37 57 38 58
rect 38 57 39 58
rect 249 57 250 58
rect 250 57 251 58
rect 251 57 252 58
rect 252 57 253 58
rect 253 57 254 58
rect 254 57 255 58
rect 255 57 256 58
rect 256 57 257 58
rect 257 57 258 58
rect 283 57 284 58
rect 284 57 285 58
rect 285 57 286 58
rect 9 56 10 57
rect 10 56 11 57
rect 11 56 12 57
rect 12 56 13 57
rect 13 56 14 57
rect 14 56 15 57
rect 15 56 16 57
rect 33 56 34 57
rect 34 56 35 57
rect 35 56 36 57
rect 36 56 37 57
rect 37 56 38 57
rect 38 56 39 57
rect 39 56 40 57
rect 249 56 250 57
rect 250 56 251 57
rect 251 56 252 57
rect 252 56 253 57
rect 253 56 254 57
rect 254 56 255 57
rect 255 56 256 57
rect 256 56 257 57
rect 282 56 283 57
rect 283 56 284 57
rect 284 56 285 57
rect 285 56 286 57
rect 9 55 10 56
rect 10 55 11 56
rect 11 55 12 56
rect 12 55 13 56
rect 13 55 14 56
rect 14 55 15 56
rect 15 55 16 56
rect 33 55 34 56
rect 34 55 35 56
rect 35 55 36 56
rect 36 55 37 56
rect 37 55 38 56
rect 38 55 39 56
rect 39 55 40 56
rect 40 55 41 56
rect 250 55 251 56
rect 251 55 252 56
rect 252 55 253 56
rect 253 55 254 56
rect 254 55 255 56
rect 255 55 256 56
rect 256 55 257 56
rect 257 55 258 56
rect 282 55 283 56
rect 283 55 284 56
rect 284 55 285 56
rect 9 54 10 55
rect 10 54 11 55
rect 11 54 12 55
rect 12 54 13 55
rect 13 54 14 55
rect 14 54 15 55
rect 15 54 16 55
rect 34 54 35 55
rect 35 54 36 55
rect 36 54 37 55
rect 37 54 38 55
rect 38 54 39 55
rect 39 54 40 55
rect 40 54 41 55
rect 250 54 251 55
rect 251 54 252 55
rect 252 54 253 55
rect 253 54 254 55
rect 254 54 255 55
rect 255 54 256 55
rect 256 54 257 55
rect 257 54 258 55
rect 281 54 282 55
rect 282 54 283 55
rect 283 54 284 55
rect 9 53 10 54
rect 10 53 11 54
rect 11 53 12 54
rect 12 53 13 54
rect 13 53 14 54
rect 14 53 15 54
rect 15 53 16 54
rect 34 53 35 54
rect 35 53 36 54
rect 36 53 37 54
rect 37 53 38 54
rect 38 53 39 54
rect 39 53 40 54
rect 40 53 41 54
rect 251 53 252 54
rect 252 53 253 54
rect 253 53 254 54
rect 254 53 255 54
rect 255 53 256 54
rect 256 53 257 54
rect 257 53 258 54
rect 258 53 259 54
rect 281 53 282 54
rect 282 53 283 54
rect 283 53 284 54
rect 9 52 10 53
rect 10 52 11 53
rect 11 52 12 53
rect 12 52 13 53
rect 13 52 14 53
rect 14 52 15 53
rect 15 52 16 53
rect 34 52 35 53
rect 35 52 36 53
rect 36 52 37 53
rect 37 52 38 53
rect 38 52 39 53
rect 39 52 40 53
rect 40 52 41 53
rect 251 52 252 53
rect 252 52 253 53
rect 253 52 254 53
rect 254 52 255 53
rect 255 52 256 53
rect 256 52 257 53
rect 257 52 258 53
rect 258 52 259 53
rect 280 52 281 53
rect 281 52 282 53
rect 282 52 283 53
rect 283 52 284 53
rect 9 51 10 52
rect 10 51 11 52
rect 11 51 12 52
rect 12 51 13 52
rect 13 51 14 52
rect 14 51 15 52
rect 15 51 16 52
rect 34 51 35 52
rect 35 51 36 52
rect 36 51 37 52
rect 37 51 38 52
rect 38 51 39 52
rect 39 51 40 52
rect 40 51 41 52
rect 252 51 253 52
rect 253 51 254 52
rect 254 51 255 52
rect 255 51 256 52
rect 256 51 257 52
rect 257 51 258 52
rect 258 51 259 52
rect 259 51 260 52
rect 280 51 281 52
rect 281 51 282 52
rect 282 51 283 52
rect 9 50 10 51
rect 10 50 11 51
rect 11 50 12 51
rect 12 50 13 51
rect 13 50 14 51
rect 14 50 15 51
rect 15 50 16 51
rect 34 50 35 51
rect 35 50 36 51
rect 36 50 37 51
rect 37 50 38 51
rect 38 50 39 51
rect 39 50 40 51
rect 40 50 41 51
rect 252 50 253 51
rect 253 50 254 51
rect 254 50 255 51
rect 255 50 256 51
rect 256 50 257 51
rect 257 50 258 51
rect 258 50 259 51
rect 259 50 260 51
rect 280 50 281 51
rect 281 50 282 51
rect 282 50 283 51
rect 283 50 284 51
rect 9 49 10 50
rect 10 49 11 50
rect 11 49 12 50
rect 12 49 13 50
rect 13 49 14 50
rect 14 49 15 50
rect 15 49 16 50
rect 34 49 35 50
rect 35 49 36 50
rect 36 49 37 50
rect 37 49 38 50
rect 38 49 39 50
rect 39 49 40 50
rect 40 49 41 50
rect 253 49 254 50
rect 254 49 255 50
rect 255 49 256 50
rect 256 49 257 50
rect 257 49 258 50
rect 258 49 259 50
rect 259 49 260 50
rect 279 49 280 50
rect 280 49 281 50
rect 281 49 282 50
rect 282 49 283 50
rect 9 48 10 49
rect 10 48 11 49
rect 11 48 12 49
rect 12 48 13 49
rect 13 48 14 49
rect 14 48 15 49
rect 15 48 16 49
rect 33 48 34 49
rect 34 48 35 49
rect 35 48 36 49
rect 36 48 37 49
rect 37 48 38 49
rect 38 48 39 49
rect 39 48 40 49
rect 40 48 41 49
rect 50 48 51 49
rect 51 48 52 49
rect 53 48 54 49
rect 55 48 56 49
rect 56 48 57 49
rect 58 48 59 49
rect 60 48 61 49
rect 69 48 70 49
rect 70 48 71 49
rect 72 48 73 49
rect 74 48 75 49
rect 75 48 76 49
rect 77 48 78 49
rect 79 48 80 49
rect 98 48 99 49
rect 99 48 100 49
rect 100 48 101 49
rect 101 48 102 49
rect 102 48 103 49
rect 103 48 104 49
rect 104 48 105 49
rect 105 48 106 49
rect 106 48 107 49
rect 108 48 109 49
rect 134 48 135 49
rect 135 48 136 49
rect 136 48 137 49
rect 137 48 138 49
rect 138 48 139 49
rect 139 48 140 49
rect 140 48 141 49
rect 141 48 142 49
rect 142 48 143 49
rect 144 48 145 49
rect 155 48 156 49
rect 157 48 158 49
rect 159 48 160 49
rect 160 48 161 49
rect 162 48 163 49
rect 164 48 165 49
rect 165 48 166 49
rect 167 48 168 49
rect 169 48 170 49
rect 179 48 180 49
rect 181 48 182 49
rect 183 48 184 49
rect 184 48 185 49
rect 186 48 187 49
rect 188 48 189 49
rect 202 48 203 49
rect 204 48 205 49
rect 205 48 206 49
rect 206 48 207 49
rect 207 48 208 49
rect 208 48 209 49
rect 209 48 210 49
rect 210 48 211 49
rect 211 48 212 49
rect 213 48 214 49
rect 253 48 254 49
rect 254 48 255 49
rect 255 48 256 49
rect 256 48 257 49
rect 257 48 258 49
rect 258 48 259 49
rect 259 48 260 49
rect 260 48 261 49
rect 278 48 279 49
rect 279 48 280 49
rect 280 48 281 49
rect 281 48 282 49
rect 282 48 283 49
rect 9 47 10 48
rect 10 47 11 48
rect 11 47 12 48
rect 12 47 13 48
rect 13 47 14 48
rect 14 47 15 48
rect 15 47 16 48
rect 33 47 34 48
rect 34 47 35 48
rect 35 47 36 48
rect 36 47 37 48
rect 37 47 38 48
rect 38 47 39 48
rect 39 47 40 48
rect 53 47 54 48
rect 54 47 55 48
rect 55 47 56 48
rect 56 47 57 48
rect 57 47 58 48
rect 58 47 59 48
rect 59 47 60 48
rect 60 47 61 48
rect 71 47 72 48
rect 72 47 73 48
rect 73 47 74 48
rect 74 47 75 48
rect 75 47 76 48
rect 76 47 77 48
rect 77 47 78 48
rect 78 47 79 48
rect 79 47 80 48
rect 95 47 96 48
rect 96 47 97 48
rect 97 47 98 48
rect 98 47 99 48
rect 104 47 105 48
rect 105 47 106 48
rect 106 47 107 48
rect 107 47 108 48
rect 108 47 109 48
rect 109 47 110 48
rect 110 47 111 48
rect 131 47 132 48
rect 132 47 133 48
rect 133 47 134 48
rect 134 47 135 48
rect 135 47 136 48
rect 136 47 137 48
rect 137 47 138 48
rect 138 47 139 48
rect 139 47 140 48
rect 140 47 141 48
rect 141 47 142 48
rect 142 47 143 48
rect 143 47 144 48
rect 144 47 145 48
rect 145 47 146 48
rect 158 47 159 48
rect 159 47 160 48
rect 160 47 161 48
rect 161 47 162 48
rect 162 47 163 48
rect 163 47 164 48
rect 164 47 165 48
rect 165 47 166 48
rect 166 47 167 48
rect 167 47 168 48
rect 168 47 169 48
rect 169 47 170 48
rect 179 47 180 48
rect 180 47 181 48
rect 181 47 182 48
rect 182 47 183 48
rect 183 47 184 48
rect 184 47 185 48
rect 185 47 186 48
rect 186 47 187 48
rect 200 47 201 48
rect 201 47 202 48
rect 202 47 203 48
rect 203 47 204 48
rect 204 47 205 48
rect 205 47 206 48
rect 206 47 207 48
rect 207 47 208 48
rect 208 47 209 48
rect 209 47 210 48
rect 210 47 211 48
rect 211 47 212 48
rect 212 47 213 48
rect 213 47 214 48
rect 214 47 215 48
rect 254 47 255 48
rect 255 47 256 48
rect 256 47 257 48
rect 257 47 258 48
rect 258 47 259 48
rect 259 47 260 48
rect 260 47 261 48
rect 261 47 262 48
rect 278 47 279 48
rect 279 47 280 48
rect 280 47 281 48
rect 281 47 282 48
rect 9 46 10 47
rect 10 46 11 47
rect 11 46 12 47
rect 12 46 13 47
rect 13 46 14 47
rect 14 46 15 47
rect 15 46 16 47
rect 32 46 33 47
rect 33 46 34 47
rect 34 46 35 47
rect 35 46 36 47
rect 36 46 37 47
rect 37 46 38 47
rect 38 46 39 47
rect 39 46 40 47
rect 54 46 55 47
rect 55 46 56 47
rect 56 46 57 47
rect 57 46 58 47
rect 58 46 59 47
rect 59 46 60 47
rect 60 46 61 47
rect 72 46 73 47
rect 73 46 74 47
rect 74 46 75 47
rect 75 46 76 47
rect 76 46 77 47
rect 77 46 78 47
rect 78 46 79 47
rect 79 46 80 47
rect 94 46 95 47
rect 95 46 96 47
rect 96 46 97 47
rect 97 46 98 47
rect 105 46 106 47
rect 106 46 107 47
rect 107 46 108 47
rect 108 46 109 47
rect 109 46 110 47
rect 110 46 111 47
rect 111 46 112 47
rect 112 46 113 47
rect 113 46 114 47
rect 114 46 115 47
rect 115 46 116 47
rect 116 46 117 47
rect 117 46 118 47
rect 118 46 119 47
rect 130 46 131 47
rect 131 46 132 47
rect 132 46 133 47
rect 133 46 134 47
rect 140 46 141 47
rect 141 46 142 47
rect 142 46 143 47
rect 143 46 144 47
rect 144 46 145 47
rect 145 46 146 47
rect 146 46 147 47
rect 147 46 148 47
rect 159 46 160 47
rect 160 46 161 47
rect 161 46 162 47
rect 162 46 163 47
rect 163 46 164 47
rect 164 46 165 47
rect 165 46 166 47
rect 182 46 183 47
rect 183 46 184 47
rect 184 46 185 47
rect 185 46 186 47
rect 186 46 187 47
rect 199 46 200 47
rect 200 46 201 47
rect 201 46 202 47
rect 202 46 203 47
rect 209 46 210 47
rect 210 46 211 47
rect 211 46 212 47
rect 212 46 213 47
rect 213 46 214 47
rect 214 46 215 47
rect 215 46 216 47
rect 216 46 217 47
rect 254 46 255 47
rect 255 46 256 47
rect 256 46 257 47
rect 257 46 258 47
rect 258 46 259 47
rect 259 46 260 47
rect 260 46 261 47
rect 261 46 262 47
rect 278 46 279 47
rect 279 46 280 47
rect 280 46 281 47
rect 281 46 282 47
rect 9 45 10 46
rect 10 45 11 46
rect 11 45 12 46
rect 12 45 13 46
rect 13 45 14 46
rect 14 45 15 46
rect 15 45 16 46
rect 31 45 32 46
rect 32 45 33 46
rect 33 45 34 46
rect 34 45 35 46
rect 35 45 36 46
rect 36 45 37 46
rect 37 45 38 46
rect 38 45 39 46
rect 54 45 55 46
rect 55 45 56 46
rect 56 45 57 46
rect 57 45 58 46
rect 58 45 59 46
rect 59 45 60 46
rect 60 45 61 46
rect 73 45 74 46
rect 74 45 75 46
rect 75 45 76 46
rect 76 45 77 46
rect 77 45 78 46
rect 78 45 79 46
rect 79 45 80 46
rect 93 45 94 46
rect 94 45 95 46
rect 95 45 96 46
rect 96 45 97 46
rect 97 45 98 46
rect 106 45 107 46
rect 107 45 108 46
rect 108 45 109 46
rect 109 45 110 46
rect 110 45 111 46
rect 111 45 112 46
rect 112 45 113 46
rect 113 45 114 46
rect 114 45 115 46
rect 115 45 116 46
rect 116 45 117 46
rect 117 45 118 46
rect 118 45 119 46
rect 129 45 130 46
rect 130 45 131 46
rect 131 45 132 46
rect 142 45 143 46
rect 143 45 144 46
rect 144 45 145 46
rect 145 45 146 46
rect 146 45 147 46
rect 147 45 148 46
rect 159 45 160 46
rect 160 45 161 46
rect 161 45 162 46
rect 162 45 163 46
rect 163 45 164 46
rect 164 45 165 46
rect 165 45 166 46
rect 182 45 183 46
rect 183 45 184 46
rect 184 45 185 46
rect 185 45 186 46
rect 198 45 199 46
rect 199 45 200 46
rect 200 45 201 46
rect 211 45 212 46
rect 212 45 213 46
rect 213 45 214 46
rect 214 45 215 46
rect 215 45 216 46
rect 216 45 217 46
rect 255 45 256 46
rect 256 45 257 46
rect 257 45 258 46
rect 258 45 259 46
rect 259 45 260 46
rect 260 45 261 46
rect 261 45 262 46
rect 262 45 263 46
rect 277 45 278 46
rect 278 45 279 46
rect 279 45 280 46
rect 280 45 281 46
rect 9 44 10 45
rect 10 44 11 45
rect 11 44 12 45
rect 12 44 13 45
rect 13 44 14 45
rect 14 44 15 45
rect 15 44 16 45
rect 30 44 31 45
rect 31 44 32 45
rect 32 44 33 45
rect 33 44 34 45
rect 34 44 35 45
rect 35 44 36 45
rect 36 44 37 45
rect 37 44 38 45
rect 55 44 56 45
rect 56 44 57 45
rect 57 44 58 45
rect 58 44 59 45
rect 59 44 60 45
rect 60 44 61 45
rect 73 44 74 45
rect 74 44 75 45
rect 75 44 76 45
rect 76 44 77 45
rect 77 44 78 45
rect 78 44 79 45
rect 79 44 80 45
rect 92 44 93 45
rect 93 44 94 45
rect 94 44 95 45
rect 95 44 96 45
rect 96 44 97 45
rect 107 44 108 45
rect 108 44 109 45
rect 109 44 110 45
rect 110 44 111 45
rect 111 44 112 45
rect 112 44 113 45
rect 113 44 114 45
rect 114 44 115 45
rect 115 44 116 45
rect 116 44 117 45
rect 117 44 118 45
rect 118 44 119 45
rect 128 44 129 45
rect 129 44 130 45
rect 130 44 131 45
rect 142 44 143 45
rect 143 44 144 45
rect 144 44 145 45
rect 145 44 146 45
rect 146 44 147 45
rect 147 44 148 45
rect 148 44 149 45
rect 160 44 161 45
rect 161 44 162 45
rect 162 44 163 45
rect 163 44 164 45
rect 164 44 165 45
rect 165 44 166 45
rect 182 44 183 45
rect 183 44 184 45
rect 184 44 185 45
rect 185 44 186 45
rect 197 44 198 45
rect 198 44 199 45
rect 199 44 200 45
rect 212 44 213 45
rect 213 44 214 45
rect 214 44 215 45
rect 215 44 216 45
rect 216 44 217 45
rect 217 44 218 45
rect 255 44 256 45
rect 256 44 257 45
rect 257 44 258 45
rect 258 44 259 45
rect 259 44 260 45
rect 260 44 261 45
rect 261 44 262 45
rect 262 44 263 45
rect 277 44 278 45
rect 278 44 279 45
rect 279 44 280 45
rect 280 44 281 45
rect 9 43 10 44
rect 10 43 11 44
rect 11 43 12 44
rect 12 43 13 44
rect 13 43 14 44
rect 14 43 15 44
rect 15 43 16 44
rect 28 43 29 44
rect 29 43 30 44
rect 30 43 31 44
rect 31 43 32 44
rect 32 43 33 44
rect 33 43 34 44
rect 34 43 35 44
rect 35 43 36 44
rect 36 43 37 44
rect 54 43 55 44
rect 55 43 56 44
rect 56 43 57 44
rect 57 43 58 44
rect 58 43 59 44
rect 59 43 60 44
rect 60 43 61 44
rect 73 43 74 44
rect 74 43 75 44
rect 75 43 76 44
rect 76 43 77 44
rect 77 43 78 44
rect 78 43 79 44
rect 79 43 80 44
rect 91 43 92 44
rect 92 43 93 44
rect 93 43 94 44
rect 94 43 95 44
rect 95 43 96 44
rect 96 43 97 44
rect 107 43 108 44
rect 108 43 109 44
rect 109 43 110 44
rect 110 43 111 44
rect 111 43 112 44
rect 112 43 113 44
rect 113 43 114 44
rect 127 43 128 44
rect 128 43 129 44
rect 129 43 130 44
rect 130 43 131 44
rect 143 43 144 44
rect 144 43 145 44
rect 145 43 146 44
rect 146 43 147 44
rect 147 43 148 44
rect 148 43 149 44
rect 149 43 150 44
rect 160 43 161 44
rect 161 43 162 44
rect 162 43 163 44
rect 163 43 164 44
rect 164 43 165 44
rect 165 43 166 44
rect 166 43 167 44
rect 182 43 183 44
rect 183 43 184 44
rect 184 43 185 44
rect 196 43 197 44
rect 197 43 198 44
rect 198 43 199 44
rect 199 43 200 44
rect 212 43 213 44
rect 213 43 214 44
rect 214 43 215 44
rect 215 43 216 44
rect 216 43 217 44
rect 217 43 218 44
rect 218 43 219 44
rect 256 43 257 44
rect 257 43 258 44
rect 258 43 259 44
rect 259 43 260 44
rect 260 43 261 44
rect 261 43 262 44
rect 262 43 263 44
rect 263 43 264 44
rect 276 43 277 44
rect 277 43 278 44
rect 278 43 279 44
rect 279 43 280 44
rect 280 43 281 44
rect 9 42 10 43
rect 10 42 11 43
rect 11 42 12 43
rect 12 42 13 43
rect 13 42 14 43
rect 14 42 15 43
rect 15 42 16 43
rect 16 42 17 43
rect 17 42 18 43
rect 18 42 19 43
rect 19 42 20 43
rect 20 42 21 43
rect 21 42 22 43
rect 22 42 23 43
rect 23 42 24 43
rect 24 42 25 43
rect 25 42 26 43
rect 26 42 27 43
rect 27 42 28 43
rect 28 42 29 43
rect 29 42 30 43
rect 30 42 31 43
rect 31 42 32 43
rect 32 42 33 43
rect 33 42 34 43
rect 34 42 35 43
rect 35 42 36 43
rect 55 42 56 43
rect 56 42 57 43
rect 57 42 58 43
rect 58 42 59 43
rect 59 42 60 43
rect 60 42 61 43
rect 73 42 74 43
rect 74 42 75 43
rect 75 42 76 43
rect 76 42 77 43
rect 77 42 78 43
rect 78 42 79 43
rect 79 42 80 43
rect 91 42 92 43
rect 92 42 93 43
rect 93 42 94 43
rect 94 42 95 43
rect 95 42 96 43
rect 96 42 97 43
rect 108 42 109 43
rect 109 42 110 43
rect 110 42 111 43
rect 111 42 112 43
rect 112 42 113 43
rect 113 42 114 43
rect 126 42 127 43
rect 127 42 128 43
rect 128 42 129 43
rect 129 42 130 43
rect 143 42 144 43
rect 144 42 145 43
rect 145 42 146 43
rect 146 42 147 43
rect 147 42 148 43
rect 148 42 149 43
rect 149 42 150 43
rect 160 42 161 43
rect 161 42 162 43
rect 162 42 163 43
rect 163 42 164 43
rect 164 42 165 43
rect 165 42 166 43
rect 166 42 167 43
rect 181 42 182 43
rect 182 42 183 43
rect 183 42 184 43
rect 184 42 185 43
rect 195 42 196 43
rect 196 42 197 43
rect 197 42 198 43
rect 198 42 199 43
rect 213 42 214 43
rect 214 42 215 43
rect 215 42 216 43
rect 216 42 217 43
rect 217 42 218 43
rect 218 42 219 43
rect 256 42 257 43
rect 257 42 258 43
rect 258 42 259 43
rect 259 42 260 43
rect 260 42 261 43
rect 261 42 262 43
rect 262 42 263 43
rect 263 42 264 43
rect 276 42 277 43
rect 277 42 278 43
rect 278 42 279 43
rect 279 42 280 43
rect 9 41 10 42
rect 10 41 11 42
rect 11 41 12 42
rect 12 41 13 42
rect 13 41 14 42
rect 14 41 15 42
rect 15 41 16 42
rect 16 41 17 42
rect 17 41 18 42
rect 18 41 19 42
rect 19 41 20 42
rect 20 41 21 42
rect 21 41 22 42
rect 22 41 23 42
rect 23 41 24 42
rect 24 41 25 42
rect 25 41 26 42
rect 26 41 27 42
rect 27 41 28 42
rect 28 41 29 42
rect 29 41 30 42
rect 30 41 31 42
rect 31 41 32 42
rect 32 41 33 42
rect 54 41 55 42
rect 55 41 56 42
rect 56 41 57 42
rect 57 41 58 42
rect 58 41 59 42
rect 59 41 60 42
rect 60 41 61 42
rect 73 41 74 42
rect 74 41 75 42
rect 75 41 76 42
rect 76 41 77 42
rect 77 41 78 42
rect 78 41 79 42
rect 79 41 80 42
rect 90 41 91 42
rect 91 41 92 42
rect 92 41 93 42
rect 93 41 94 42
rect 94 41 95 42
rect 95 41 96 42
rect 107 41 108 42
rect 108 41 109 42
rect 109 41 110 42
rect 110 41 111 42
rect 111 41 112 42
rect 112 41 113 42
rect 113 41 114 42
rect 126 41 127 42
rect 127 41 128 42
rect 128 41 129 42
rect 129 41 130 42
rect 143 41 144 42
rect 144 41 145 42
rect 145 41 146 42
rect 146 41 147 42
rect 147 41 148 42
rect 148 41 149 42
rect 149 41 150 42
rect 150 41 151 42
rect 161 41 162 42
rect 162 41 163 42
rect 163 41 164 42
rect 164 41 165 42
rect 165 41 166 42
rect 166 41 167 42
rect 167 41 168 42
rect 181 41 182 42
rect 182 41 183 42
rect 183 41 184 42
rect 196 41 197 42
rect 197 41 198 42
rect 198 41 199 42
rect 213 41 214 42
rect 214 41 215 42
rect 215 41 216 42
rect 216 41 217 42
rect 217 41 218 42
rect 218 41 219 42
rect 219 41 220 42
rect 257 41 258 42
rect 258 41 259 42
rect 259 41 260 42
rect 260 41 261 42
rect 261 41 262 42
rect 262 41 263 42
rect 263 41 264 42
rect 276 41 277 42
rect 277 41 278 42
rect 278 41 279 42
rect 279 41 280 42
rect 9 40 10 41
rect 10 40 11 41
rect 11 40 12 41
rect 12 40 13 41
rect 13 40 14 41
rect 14 40 15 41
rect 15 40 16 41
rect 16 40 17 41
rect 17 40 18 41
rect 18 40 19 41
rect 19 40 20 41
rect 20 40 21 41
rect 21 40 22 41
rect 22 40 23 41
rect 23 40 24 41
rect 24 40 25 41
rect 25 40 26 41
rect 26 40 27 41
rect 27 40 28 41
rect 28 40 29 41
rect 29 40 30 41
rect 30 40 31 41
rect 31 40 32 41
rect 32 40 33 41
rect 33 40 34 41
rect 34 40 35 41
rect 54 40 55 41
rect 55 40 56 41
rect 56 40 57 41
rect 57 40 58 41
rect 58 40 59 41
rect 59 40 60 41
rect 60 40 61 41
rect 73 40 74 41
rect 74 40 75 41
rect 75 40 76 41
rect 76 40 77 41
rect 77 40 78 41
rect 78 40 79 41
rect 79 40 80 41
rect 90 40 91 41
rect 91 40 92 41
rect 92 40 93 41
rect 93 40 94 41
rect 94 40 95 41
rect 95 40 96 41
rect 108 40 109 41
rect 109 40 110 41
rect 110 40 111 41
rect 111 40 112 41
rect 112 40 113 41
rect 113 40 114 41
rect 114 40 115 41
rect 125 40 126 41
rect 126 40 127 41
rect 127 40 128 41
rect 128 40 129 41
rect 129 40 130 41
rect 143 40 144 41
rect 144 40 145 41
rect 145 40 146 41
rect 146 40 147 41
rect 147 40 148 41
rect 148 40 149 41
rect 149 40 150 41
rect 150 40 151 41
rect 161 40 162 41
rect 162 40 163 41
rect 163 40 164 41
rect 164 40 165 41
rect 165 40 166 41
rect 166 40 167 41
rect 167 40 168 41
rect 180 40 181 41
rect 181 40 182 41
rect 182 40 183 41
rect 183 40 184 41
rect 195 40 196 41
rect 196 40 197 41
rect 197 40 198 41
rect 198 40 199 41
rect 213 40 214 41
rect 214 40 215 41
rect 215 40 216 41
rect 216 40 217 41
rect 217 40 218 41
rect 218 40 219 41
rect 219 40 220 41
rect 257 40 258 41
rect 258 40 259 41
rect 259 40 260 41
rect 260 40 261 41
rect 261 40 262 41
rect 262 40 263 41
rect 263 40 264 41
rect 264 40 265 41
rect 275 40 276 41
rect 276 40 277 41
rect 277 40 278 41
rect 278 40 279 41
rect 9 39 10 40
rect 10 39 11 40
rect 11 39 12 40
rect 12 39 13 40
rect 13 39 14 40
rect 14 39 15 40
rect 15 39 16 40
rect 27 39 28 40
rect 28 39 29 40
rect 29 39 30 40
rect 30 39 31 40
rect 31 39 32 40
rect 32 39 33 40
rect 33 39 34 40
rect 34 39 35 40
rect 35 39 36 40
rect 36 39 37 40
rect 37 39 38 40
rect 55 39 56 40
rect 56 39 57 40
rect 57 39 58 40
rect 58 39 59 40
rect 59 39 60 40
rect 60 39 61 40
rect 73 39 74 40
rect 74 39 75 40
rect 75 39 76 40
rect 76 39 77 40
rect 77 39 78 40
rect 78 39 79 40
rect 79 39 80 40
rect 89 39 90 40
rect 90 39 91 40
rect 91 39 92 40
rect 92 39 93 40
rect 93 39 94 40
rect 94 39 95 40
rect 95 39 96 40
rect 108 39 109 40
rect 109 39 110 40
rect 110 39 111 40
rect 111 39 112 40
rect 112 39 113 40
rect 113 39 114 40
rect 114 39 115 40
rect 124 39 125 40
rect 125 39 126 40
rect 126 39 127 40
rect 127 39 128 40
rect 128 39 129 40
rect 144 39 145 40
rect 145 39 146 40
rect 146 39 147 40
rect 147 39 148 40
rect 148 39 149 40
rect 149 39 150 40
rect 150 39 151 40
rect 162 39 163 40
rect 163 39 164 40
rect 164 39 165 40
rect 165 39 166 40
rect 166 39 167 40
rect 167 39 168 40
rect 168 39 169 40
rect 180 39 181 40
rect 181 39 182 40
rect 182 39 183 40
rect 194 39 195 40
rect 195 39 196 40
rect 196 39 197 40
rect 197 39 198 40
rect 213 39 214 40
rect 214 39 215 40
rect 215 39 216 40
rect 216 39 217 40
rect 217 39 218 40
rect 218 39 219 40
rect 219 39 220 40
rect 258 39 259 40
rect 259 39 260 40
rect 260 39 261 40
rect 261 39 262 40
rect 262 39 263 40
rect 263 39 264 40
rect 264 39 265 40
rect 265 39 266 40
rect 274 39 275 40
rect 275 39 276 40
rect 276 39 277 40
rect 277 39 278 40
rect 278 39 279 40
rect 9 38 10 39
rect 10 38 11 39
rect 11 38 12 39
rect 12 38 13 39
rect 13 38 14 39
rect 14 38 15 39
rect 15 38 16 39
rect 30 38 31 39
rect 31 38 32 39
rect 32 38 33 39
rect 33 38 34 39
rect 34 38 35 39
rect 35 38 36 39
rect 36 38 37 39
rect 37 38 38 39
rect 38 38 39 39
rect 54 38 55 39
rect 55 38 56 39
rect 56 38 57 39
rect 57 38 58 39
rect 58 38 59 39
rect 59 38 60 39
rect 60 38 61 39
rect 73 38 74 39
rect 74 38 75 39
rect 75 38 76 39
rect 76 38 77 39
rect 77 38 78 39
rect 78 38 79 39
rect 79 38 80 39
rect 90 38 91 39
rect 91 38 92 39
rect 92 38 93 39
rect 93 38 94 39
rect 94 38 95 39
rect 95 38 96 39
rect 108 38 109 39
rect 109 38 110 39
rect 110 38 111 39
rect 111 38 112 39
rect 112 38 113 39
rect 113 38 114 39
rect 114 38 115 39
rect 125 38 126 39
rect 126 38 127 39
rect 127 38 128 39
rect 128 38 129 39
rect 129 38 130 39
rect 130 38 131 39
rect 131 38 132 39
rect 132 38 133 39
rect 133 38 134 39
rect 134 38 135 39
rect 135 38 136 39
rect 136 38 137 39
rect 137 38 138 39
rect 138 38 139 39
rect 139 38 140 39
rect 140 38 141 39
rect 141 38 142 39
rect 142 38 143 39
rect 143 38 144 39
rect 144 38 145 39
rect 145 38 146 39
rect 146 38 147 39
rect 147 38 148 39
rect 148 38 149 39
rect 149 38 150 39
rect 150 38 151 39
rect 151 38 152 39
rect 162 38 163 39
rect 163 38 164 39
rect 164 38 165 39
rect 165 38 166 39
rect 166 38 167 39
rect 167 38 168 39
rect 180 38 181 39
rect 181 38 182 39
rect 182 38 183 39
rect 194 38 195 39
rect 195 38 196 39
rect 196 38 197 39
rect 197 38 198 39
rect 198 38 199 39
rect 199 38 200 39
rect 200 38 201 39
rect 201 38 202 39
rect 202 38 203 39
rect 203 38 204 39
rect 204 38 205 39
rect 205 38 206 39
rect 206 38 207 39
rect 207 38 208 39
rect 208 38 209 39
rect 209 38 210 39
rect 210 38 211 39
rect 211 38 212 39
rect 212 38 213 39
rect 213 38 214 39
rect 214 38 215 39
rect 215 38 216 39
rect 216 38 217 39
rect 217 38 218 39
rect 218 38 219 39
rect 219 38 220 39
rect 220 38 221 39
rect 257 38 258 39
rect 258 38 259 39
rect 259 38 260 39
rect 260 38 261 39
rect 261 38 262 39
rect 262 38 263 39
rect 263 38 264 39
rect 264 38 265 39
rect 275 38 276 39
rect 276 38 277 39
rect 277 38 278 39
rect 9 37 10 38
rect 10 37 11 38
rect 11 37 12 38
rect 12 37 13 38
rect 13 37 14 38
rect 14 37 15 38
rect 15 37 16 38
rect 31 37 32 38
rect 32 37 33 38
rect 33 37 34 38
rect 34 37 35 38
rect 35 37 36 38
rect 36 37 37 38
rect 37 37 38 38
rect 38 37 39 38
rect 39 37 40 38
rect 55 37 56 38
rect 56 37 57 38
rect 57 37 58 38
rect 58 37 59 38
rect 59 37 60 38
rect 60 37 61 38
rect 73 37 74 38
rect 74 37 75 38
rect 75 37 76 38
rect 76 37 77 38
rect 77 37 78 38
rect 78 37 79 38
rect 79 37 80 38
rect 89 37 90 38
rect 90 37 91 38
rect 91 37 92 38
rect 92 37 93 38
rect 93 37 94 38
rect 94 37 95 38
rect 95 37 96 38
rect 96 37 97 38
rect 108 37 109 38
rect 109 37 110 38
rect 110 37 111 38
rect 111 37 112 38
rect 112 37 113 38
rect 113 37 114 38
rect 114 37 115 38
rect 124 37 125 38
rect 125 37 126 38
rect 126 37 127 38
rect 127 37 128 38
rect 128 37 129 38
rect 129 37 130 38
rect 130 37 131 38
rect 131 37 132 38
rect 132 37 133 38
rect 133 37 134 38
rect 134 37 135 38
rect 135 37 136 38
rect 136 37 137 38
rect 137 37 138 38
rect 138 37 139 38
rect 139 37 140 38
rect 140 37 141 38
rect 141 37 142 38
rect 142 37 143 38
rect 143 37 144 38
rect 144 37 145 38
rect 145 37 146 38
rect 146 37 147 38
rect 147 37 148 38
rect 148 37 149 38
rect 149 37 150 38
rect 150 37 151 38
rect 163 37 164 38
rect 164 37 165 38
rect 165 37 166 38
rect 166 37 167 38
rect 167 37 168 38
rect 168 37 169 38
rect 179 37 180 38
rect 180 37 181 38
rect 181 37 182 38
rect 182 37 183 38
rect 194 37 195 38
rect 195 37 196 38
rect 196 37 197 38
rect 197 37 198 38
rect 198 37 199 38
rect 199 37 200 38
rect 200 37 201 38
rect 201 37 202 38
rect 202 37 203 38
rect 203 37 204 38
rect 204 37 205 38
rect 205 37 206 38
rect 206 37 207 38
rect 207 37 208 38
rect 208 37 209 38
rect 209 37 210 38
rect 210 37 211 38
rect 211 37 212 38
rect 212 37 213 38
rect 213 37 214 38
rect 214 37 215 38
rect 215 37 216 38
rect 216 37 217 38
rect 217 37 218 38
rect 218 37 219 38
rect 219 37 220 38
rect 220 37 221 38
rect 258 37 259 38
rect 259 37 260 38
rect 260 37 261 38
rect 261 37 262 38
rect 262 37 263 38
rect 263 37 264 38
rect 264 37 265 38
rect 265 37 266 38
rect 274 37 275 38
rect 275 37 276 38
rect 276 37 277 38
rect 277 37 278 38
rect 9 36 10 37
rect 10 36 11 37
rect 11 36 12 37
rect 12 36 13 37
rect 13 36 14 37
rect 14 36 15 37
rect 15 36 16 37
rect 33 36 34 37
rect 34 36 35 37
rect 35 36 36 37
rect 36 36 37 37
rect 37 36 38 37
rect 38 36 39 37
rect 39 36 40 37
rect 40 36 41 37
rect 54 36 55 37
rect 55 36 56 37
rect 56 36 57 37
rect 57 36 58 37
rect 58 36 59 37
rect 59 36 60 37
rect 60 36 61 37
rect 73 36 74 37
rect 74 36 75 37
rect 75 36 76 37
rect 76 36 77 37
rect 77 36 78 37
rect 78 36 79 37
rect 79 36 80 37
rect 90 36 91 37
rect 91 36 92 37
rect 92 36 93 37
rect 93 36 94 37
rect 94 36 95 37
rect 95 36 96 37
rect 96 36 97 37
rect 108 36 109 37
rect 109 36 110 37
rect 110 36 111 37
rect 111 36 112 37
rect 112 36 113 37
rect 113 36 114 37
rect 114 36 115 37
rect 125 36 126 37
rect 126 36 127 37
rect 127 36 128 37
rect 128 36 129 37
rect 163 36 164 37
rect 164 36 165 37
rect 165 36 166 37
rect 166 36 167 37
rect 167 36 168 37
rect 168 36 169 37
rect 179 36 180 37
rect 180 36 181 37
rect 181 36 182 37
rect 194 36 195 37
rect 195 36 196 37
rect 196 36 197 37
rect 197 36 198 37
rect 258 36 259 37
rect 259 36 260 37
rect 260 36 261 37
rect 261 36 262 37
rect 262 36 263 37
rect 263 36 264 37
rect 264 36 265 37
rect 265 36 266 37
rect 274 36 275 37
rect 275 36 276 37
rect 276 36 277 37
rect 9 35 10 36
rect 10 35 11 36
rect 11 35 12 36
rect 12 35 13 36
rect 13 35 14 36
rect 14 35 15 36
rect 15 35 16 36
rect 34 35 35 36
rect 35 35 36 36
rect 36 35 37 36
rect 37 35 38 36
rect 38 35 39 36
rect 39 35 40 36
rect 40 35 41 36
rect 41 35 42 36
rect 54 35 55 36
rect 55 35 56 36
rect 56 35 57 36
rect 57 35 58 36
rect 58 35 59 36
rect 59 35 60 36
rect 60 35 61 36
rect 73 35 74 36
rect 74 35 75 36
rect 75 35 76 36
rect 76 35 77 36
rect 77 35 78 36
rect 78 35 79 36
rect 79 35 80 36
rect 90 35 91 36
rect 91 35 92 36
rect 92 35 93 36
rect 93 35 94 36
rect 94 35 95 36
rect 95 35 96 36
rect 96 35 97 36
rect 108 35 109 36
rect 109 35 110 36
rect 110 35 111 36
rect 111 35 112 36
rect 112 35 113 36
rect 113 35 114 36
rect 114 35 115 36
rect 124 35 125 36
rect 125 35 126 36
rect 126 35 127 36
rect 127 35 128 36
rect 128 35 129 36
rect 163 35 164 36
rect 164 35 165 36
rect 165 35 166 36
rect 166 35 167 36
rect 167 35 168 36
rect 168 35 169 36
rect 169 35 170 36
rect 179 35 180 36
rect 180 35 181 36
rect 181 35 182 36
rect 193 35 194 36
rect 194 35 195 36
rect 195 35 196 36
rect 196 35 197 36
rect 197 35 198 36
rect 259 35 260 36
rect 260 35 261 36
rect 261 35 262 36
rect 262 35 263 36
rect 263 35 264 36
rect 264 35 265 36
rect 265 35 266 36
rect 266 35 267 36
rect 274 35 275 36
rect 275 35 276 36
rect 276 35 277 36
rect 9 34 10 35
rect 10 34 11 35
rect 11 34 12 35
rect 12 34 13 35
rect 13 34 14 35
rect 14 34 15 35
rect 15 34 16 35
rect 34 34 35 35
rect 35 34 36 35
rect 36 34 37 35
rect 37 34 38 35
rect 38 34 39 35
rect 39 34 40 35
rect 40 34 41 35
rect 41 34 42 35
rect 55 34 56 35
rect 56 34 57 35
rect 57 34 58 35
rect 58 34 59 35
rect 59 34 60 35
rect 60 34 61 35
rect 73 34 74 35
rect 74 34 75 35
rect 75 34 76 35
rect 76 34 77 35
rect 77 34 78 35
rect 78 34 79 35
rect 79 34 80 35
rect 90 34 91 35
rect 91 34 92 35
rect 92 34 93 35
rect 93 34 94 35
rect 94 34 95 35
rect 95 34 96 35
rect 96 34 97 35
rect 108 34 109 35
rect 109 34 110 35
rect 110 34 111 35
rect 111 34 112 35
rect 112 34 113 35
rect 113 34 114 35
rect 124 34 125 35
rect 125 34 126 35
rect 126 34 127 35
rect 127 34 128 35
rect 128 34 129 35
rect 164 34 165 35
rect 165 34 166 35
rect 166 34 167 35
rect 167 34 168 35
rect 168 34 169 35
rect 169 34 170 35
rect 178 34 179 35
rect 179 34 180 35
rect 180 34 181 35
rect 193 34 194 35
rect 194 34 195 35
rect 195 34 196 35
rect 196 34 197 35
rect 197 34 198 35
rect 259 34 260 35
rect 260 34 261 35
rect 261 34 262 35
rect 262 34 263 35
rect 263 34 264 35
rect 264 34 265 35
rect 265 34 266 35
rect 266 34 267 35
rect 273 34 274 35
rect 274 34 275 35
rect 275 34 276 35
rect 276 34 277 35
rect 9 33 10 34
rect 10 33 11 34
rect 11 33 12 34
rect 12 33 13 34
rect 13 33 14 34
rect 14 33 15 34
rect 15 33 16 34
rect 35 33 36 34
rect 36 33 37 34
rect 37 33 38 34
rect 38 33 39 34
rect 39 33 40 34
rect 40 33 41 34
rect 41 33 42 34
rect 54 33 55 34
rect 55 33 56 34
rect 56 33 57 34
rect 57 33 58 34
rect 58 33 59 34
rect 59 33 60 34
rect 60 33 61 34
rect 73 33 74 34
rect 74 33 75 34
rect 75 33 76 34
rect 76 33 77 34
rect 77 33 78 34
rect 78 33 79 34
rect 79 33 80 34
rect 90 33 91 34
rect 91 33 92 34
rect 92 33 93 34
rect 93 33 94 34
rect 94 33 95 34
rect 95 33 96 34
rect 96 33 97 34
rect 97 33 98 34
rect 108 33 109 34
rect 109 33 110 34
rect 110 33 111 34
rect 111 33 112 34
rect 112 33 113 34
rect 113 33 114 34
rect 124 33 125 34
rect 125 33 126 34
rect 126 33 127 34
rect 127 33 128 34
rect 128 33 129 34
rect 164 33 165 34
rect 165 33 166 34
rect 166 33 167 34
rect 167 33 168 34
rect 168 33 169 34
rect 169 33 170 34
rect 170 33 171 34
rect 178 33 179 34
rect 179 33 180 34
rect 180 33 181 34
rect 193 33 194 34
rect 194 33 195 34
rect 195 33 196 34
rect 196 33 197 34
rect 197 33 198 34
rect 260 33 261 34
rect 261 33 262 34
rect 262 33 263 34
rect 263 33 264 34
rect 264 33 265 34
rect 265 33 266 34
rect 266 33 267 34
rect 273 33 274 34
rect 274 33 275 34
rect 275 33 276 34
rect 9 32 10 33
rect 10 32 11 33
rect 11 32 12 33
rect 12 32 13 33
rect 13 32 14 33
rect 14 32 15 33
rect 15 32 16 33
rect 35 32 36 33
rect 36 32 37 33
rect 37 32 38 33
rect 38 32 39 33
rect 39 32 40 33
rect 40 32 41 33
rect 41 32 42 33
rect 42 32 43 33
rect 55 32 56 33
rect 56 32 57 33
rect 57 32 58 33
rect 58 32 59 33
rect 59 32 60 33
rect 60 32 61 33
rect 73 32 74 33
rect 74 32 75 33
rect 75 32 76 33
rect 76 32 77 33
rect 77 32 78 33
rect 78 32 79 33
rect 79 32 80 33
rect 91 32 92 33
rect 92 32 93 33
rect 93 32 94 33
rect 94 32 95 33
rect 95 32 96 33
rect 96 32 97 33
rect 97 32 98 33
rect 108 32 109 33
rect 109 32 110 33
rect 110 32 111 33
rect 111 32 112 33
rect 112 32 113 33
rect 113 32 114 33
rect 124 32 125 33
rect 125 32 126 33
rect 126 32 127 33
rect 127 32 128 33
rect 128 32 129 33
rect 165 32 166 33
rect 166 32 167 33
rect 167 32 168 33
rect 168 32 169 33
rect 169 32 170 33
rect 170 32 171 33
rect 171 32 172 33
rect 177 32 178 33
rect 178 32 179 33
rect 179 32 180 33
rect 180 32 181 33
rect 193 32 194 33
rect 194 32 195 33
rect 195 32 196 33
rect 196 32 197 33
rect 197 32 198 33
rect 260 32 261 33
rect 261 32 262 33
rect 262 32 263 33
rect 263 32 264 33
rect 264 32 265 33
rect 265 32 266 33
rect 266 32 267 33
rect 267 32 268 33
rect 272 32 273 33
rect 273 32 274 33
rect 274 32 275 33
rect 275 32 276 33
rect 9 31 10 32
rect 10 31 11 32
rect 11 31 12 32
rect 12 31 13 32
rect 13 31 14 32
rect 14 31 15 32
rect 15 31 16 32
rect 36 31 37 32
rect 37 31 38 32
rect 38 31 39 32
rect 39 31 40 32
rect 40 31 41 32
rect 41 31 42 32
rect 42 31 43 32
rect 54 31 55 32
rect 55 31 56 32
rect 56 31 57 32
rect 57 31 58 32
rect 58 31 59 32
rect 59 31 60 32
rect 60 31 61 32
rect 73 31 74 32
rect 74 31 75 32
rect 75 31 76 32
rect 76 31 77 32
rect 77 31 78 32
rect 78 31 79 32
rect 79 31 80 32
rect 92 31 93 32
rect 93 31 94 32
rect 94 31 95 32
rect 95 31 96 32
rect 96 31 97 32
rect 97 31 98 32
rect 98 31 99 32
rect 107 31 108 32
rect 108 31 109 32
rect 109 31 110 32
rect 110 31 111 32
rect 111 31 112 32
rect 124 31 125 32
rect 125 31 126 32
rect 126 31 127 32
rect 127 31 128 32
rect 128 31 129 32
rect 129 31 130 32
rect 166 31 167 32
rect 167 31 168 32
rect 168 31 169 32
rect 169 31 170 32
rect 170 31 171 32
rect 171 31 172 32
rect 178 31 179 32
rect 179 31 180 32
rect 193 31 194 32
rect 194 31 195 32
rect 195 31 196 32
rect 196 31 197 32
rect 197 31 198 32
rect 198 31 199 32
rect 261 31 262 32
rect 262 31 263 32
rect 263 31 264 32
rect 264 31 265 32
rect 265 31 266 32
rect 266 31 267 32
rect 267 31 268 32
rect 268 31 269 32
rect 272 31 273 32
rect 273 31 274 32
rect 274 31 275 32
rect 9 30 10 31
rect 10 30 11 31
rect 11 30 12 31
rect 12 30 13 31
rect 13 30 14 31
rect 14 30 15 31
rect 15 30 16 31
rect 36 30 37 31
rect 37 30 38 31
rect 38 30 39 31
rect 39 30 40 31
rect 40 30 41 31
rect 41 30 42 31
rect 42 30 43 31
rect 54 30 55 31
rect 55 30 56 31
rect 56 30 57 31
rect 57 30 58 31
rect 58 30 59 31
rect 59 30 60 31
rect 60 30 61 31
rect 73 30 74 31
rect 74 30 75 31
rect 75 30 76 31
rect 76 30 77 31
rect 77 30 78 31
rect 78 30 79 31
rect 79 30 80 31
rect 93 30 94 31
rect 94 30 95 31
rect 95 30 96 31
rect 96 30 97 31
rect 97 30 98 31
rect 98 30 99 31
rect 107 30 108 31
rect 108 30 109 31
rect 109 30 110 31
rect 110 30 111 31
rect 124 30 125 31
rect 125 30 126 31
rect 126 30 127 31
rect 127 30 128 31
rect 128 30 129 31
rect 129 30 130 31
rect 166 30 167 31
rect 167 30 168 31
rect 168 30 169 31
rect 169 30 170 31
rect 170 30 171 31
rect 171 30 172 31
rect 172 30 173 31
rect 177 30 178 31
rect 178 30 179 31
rect 179 30 180 31
rect 193 30 194 31
rect 194 30 195 31
rect 195 30 196 31
rect 196 30 197 31
rect 197 30 198 31
rect 198 30 199 31
rect 261 30 262 31
rect 262 30 263 31
rect 263 30 264 31
rect 264 30 265 31
rect 265 30 266 31
rect 266 30 267 31
rect 267 30 268 31
rect 268 30 269 31
rect 271 30 272 31
rect 272 30 273 31
rect 273 30 274 31
rect 274 30 275 31
rect 9 29 10 30
rect 10 29 11 30
rect 11 29 12 30
rect 12 29 13 30
rect 13 29 14 30
rect 14 29 15 30
rect 15 29 16 30
rect 36 29 37 30
rect 37 29 38 30
rect 38 29 39 30
rect 39 29 40 30
rect 40 29 41 30
rect 41 29 42 30
rect 42 29 43 30
rect 55 29 56 30
rect 56 29 57 30
rect 57 29 58 30
rect 58 29 59 30
rect 59 29 60 30
rect 60 29 61 30
rect 73 29 74 30
rect 74 29 75 30
rect 75 29 76 30
rect 76 29 77 30
rect 77 29 78 30
rect 78 29 79 30
rect 79 29 80 30
rect 95 29 96 30
rect 96 29 97 30
rect 97 29 98 30
rect 98 29 99 30
rect 99 29 100 30
rect 100 29 101 30
rect 106 29 107 30
rect 107 29 108 30
rect 108 29 109 30
rect 109 29 110 30
rect 124 29 125 30
rect 125 29 126 30
rect 126 29 127 30
rect 127 29 128 30
rect 128 29 129 30
rect 129 29 130 30
rect 167 29 168 30
rect 168 29 169 30
rect 169 29 170 30
rect 170 29 171 30
rect 171 29 172 30
rect 172 29 173 30
rect 177 29 178 30
rect 178 29 179 30
rect 193 29 194 30
rect 194 29 195 30
rect 195 29 196 30
rect 196 29 197 30
rect 197 29 198 30
rect 198 29 199 30
rect 262 29 263 30
rect 263 29 264 30
rect 264 29 265 30
rect 265 29 266 30
rect 266 29 267 30
rect 267 29 268 30
rect 268 29 269 30
rect 269 29 270 30
rect 271 29 272 30
rect 272 29 273 30
rect 273 29 274 30
rect 9 28 10 29
rect 10 28 11 29
rect 11 28 12 29
rect 12 28 13 29
rect 13 28 14 29
rect 14 28 15 29
rect 15 28 16 29
rect 36 28 37 29
rect 37 28 38 29
rect 38 28 39 29
rect 39 28 40 29
rect 40 28 41 29
rect 41 28 42 29
rect 42 28 43 29
rect 54 28 55 29
rect 55 28 56 29
rect 56 28 57 29
rect 57 28 58 29
rect 58 28 59 29
rect 59 28 60 29
rect 60 28 61 29
rect 73 28 74 29
rect 74 28 75 29
rect 75 28 76 29
rect 76 28 77 29
rect 77 28 78 29
rect 78 28 79 29
rect 79 28 80 29
rect 97 28 98 29
rect 98 28 99 29
rect 99 28 100 29
rect 100 28 101 29
rect 101 28 102 29
rect 102 28 103 29
rect 103 28 104 29
rect 104 28 105 29
rect 105 28 106 29
rect 106 28 107 29
rect 107 28 108 29
rect 124 28 125 29
rect 125 28 126 29
rect 126 28 127 29
rect 127 28 128 29
rect 128 28 129 29
rect 129 28 130 29
rect 167 28 168 29
rect 168 28 169 29
rect 169 28 170 29
rect 170 28 171 29
rect 171 28 172 29
rect 172 28 173 29
rect 177 28 178 29
rect 178 28 179 29
rect 193 28 194 29
rect 194 28 195 29
rect 195 28 196 29
rect 196 28 197 29
rect 197 28 198 29
rect 198 28 199 29
rect 262 28 263 29
rect 263 28 264 29
rect 264 28 265 29
rect 265 28 266 29
rect 266 28 267 29
rect 267 28 268 29
rect 268 28 269 29
rect 269 28 270 29
rect 271 28 272 29
rect 272 28 273 29
rect 273 28 274 29
rect 274 28 275 29
rect 9 27 10 28
rect 10 27 11 28
rect 11 27 12 28
rect 12 27 13 28
rect 13 27 14 28
rect 14 27 15 28
rect 15 27 16 28
rect 36 27 37 28
rect 37 27 38 28
rect 38 27 39 28
rect 39 27 40 28
rect 40 27 41 28
rect 41 27 42 28
rect 42 27 43 28
rect 55 27 56 28
rect 56 27 57 28
rect 57 27 58 28
rect 58 27 59 28
rect 59 27 60 28
rect 60 27 61 28
rect 73 27 74 28
rect 74 27 75 28
rect 75 27 76 28
rect 76 27 77 28
rect 77 27 78 28
rect 78 27 79 28
rect 79 27 80 28
rect 96 27 97 28
rect 97 27 98 28
rect 98 27 99 28
rect 99 27 100 28
rect 100 27 101 28
rect 101 27 102 28
rect 102 27 103 28
rect 103 27 104 28
rect 104 27 105 28
rect 105 27 106 28
rect 106 27 107 28
rect 124 27 125 28
rect 125 27 126 28
rect 126 27 127 28
rect 127 27 128 28
rect 128 27 129 28
rect 129 27 130 28
rect 130 27 131 28
rect 151 27 152 28
rect 168 27 169 28
rect 169 27 170 28
rect 170 27 171 28
rect 171 27 172 28
rect 172 27 173 28
rect 173 27 174 28
rect 176 27 177 28
rect 177 27 178 28
rect 193 27 194 28
rect 194 27 195 28
rect 195 27 196 28
rect 196 27 197 28
rect 197 27 198 28
rect 198 27 199 28
rect 199 27 200 28
rect 221 27 222 28
rect 263 27 264 28
rect 264 27 265 28
rect 265 27 266 28
rect 266 27 267 28
rect 267 27 268 28
rect 268 27 269 28
rect 269 27 270 28
rect 270 27 271 28
rect 271 27 272 28
rect 272 27 273 28
rect 273 27 274 28
rect 9 26 10 27
rect 10 26 11 27
rect 11 26 12 27
rect 12 26 13 27
rect 13 26 14 27
rect 14 26 15 27
rect 15 26 16 27
rect 36 26 37 27
rect 37 26 38 27
rect 38 26 39 27
rect 39 26 40 27
rect 40 26 41 27
rect 41 26 42 27
rect 42 26 43 27
rect 54 26 55 27
rect 55 26 56 27
rect 56 26 57 27
rect 57 26 58 27
rect 58 26 59 27
rect 59 26 60 27
rect 60 26 61 27
rect 73 26 74 27
rect 74 26 75 27
rect 75 26 76 27
rect 76 26 77 27
rect 77 26 78 27
rect 78 26 79 27
rect 79 26 80 27
rect 95 26 96 27
rect 96 26 97 27
rect 97 26 98 27
rect 124 26 125 27
rect 125 26 126 27
rect 126 26 127 27
rect 127 26 128 27
rect 128 26 129 27
rect 129 26 130 27
rect 130 26 131 27
rect 151 26 152 27
rect 168 26 169 27
rect 169 26 170 27
rect 170 26 171 27
rect 171 26 172 27
rect 172 26 173 27
rect 173 26 174 27
rect 176 26 177 27
rect 177 26 178 27
rect 194 26 195 27
rect 195 26 196 27
rect 196 26 197 27
rect 197 26 198 27
rect 198 26 199 27
rect 199 26 200 27
rect 220 26 221 27
rect 263 26 264 27
rect 264 26 265 27
rect 265 26 266 27
rect 266 26 267 27
rect 267 26 268 27
rect 268 26 269 27
rect 269 26 270 27
rect 270 26 271 27
rect 271 26 272 27
rect 272 26 273 27
rect 273 26 274 27
rect 9 25 10 26
rect 10 25 11 26
rect 11 25 12 26
rect 12 25 13 26
rect 13 25 14 26
rect 14 25 15 26
rect 15 25 16 26
rect 35 25 36 26
rect 36 25 37 26
rect 37 25 38 26
rect 38 25 39 26
rect 39 25 40 26
rect 40 25 41 26
rect 41 25 42 26
rect 42 25 43 26
rect 54 25 55 26
rect 55 25 56 26
rect 56 25 57 26
rect 57 25 58 26
rect 58 25 59 26
rect 59 25 60 26
rect 60 25 61 26
rect 73 25 74 26
rect 74 25 75 26
rect 75 25 76 26
rect 76 25 77 26
rect 77 25 78 26
rect 78 25 79 26
rect 79 25 80 26
rect 94 25 95 26
rect 95 25 96 26
rect 96 25 97 26
rect 125 25 126 26
rect 126 25 127 26
rect 127 25 128 26
rect 128 25 129 26
rect 129 25 130 26
rect 130 25 131 26
rect 131 25 132 26
rect 150 25 151 26
rect 168 25 169 26
rect 169 25 170 26
rect 170 25 171 26
rect 171 25 172 26
rect 172 25 173 26
rect 173 25 174 26
rect 174 25 175 26
rect 176 25 177 26
rect 177 25 178 26
rect 194 25 195 26
rect 195 25 196 26
rect 196 25 197 26
rect 197 25 198 26
rect 198 25 199 26
rect 199 25 200 26
rect 200 25 201 26
rect 219 25 220 26
rect 220 25 221 26
rect 264 25 265 26
rect 265 25 266 26
rect 266 25 267 26
rect 267 25 268 26
rect 268 25 269 26
rect 269 25 270 26
rect 270 25 271 26
rect 271 25 272 26
rect 272 25 273 26
rect 273 25 274 26
rect 9 24 10 25
rect 10 24 11 25
rect 11 24 12 25
rect 12 24 13 25
rect 13 24 14 25
rect 14 24 15 25
rect 15 24 16 25
rect 34 24 35 25
rect 35 24 36 25
rect 36 24 37 25
rect 37 24 38 25
rect 38 24 39 25
rect 39 24 40 25
rect 40 24 41 25
rect 41 24 42 25
rect 55 24 56 25
rect 56 24 57 25
rect 57 24 58 25
rect 58 24 59 25
rect 59 24 60 25
rect 60 24 61 25
rect 73 24 74 25
rect 74 24 75 25
rect 75 24 76 25
rect 76 24 77 25
rect 77 24 78 25
rect 78 24 79 25
rect 79 24 80 25
rect 92 24 93 25
rect 93 24 94 25
rect 94 24 95 25
rect 95 24 96 25
rect 125 24 126 25
rect 126 24 127 25
rect 127 24 128 25
rect 128 24 129 25
rect 129 24 130 25
rect 130 24 131 25
rect 131 24 132 25
rect 132 24 133 25
rect 148 24 149 25
rect 149 24 150 25
rect 150 24 151 25
rect 169 24 170 25
rect 170 24 171 25
rect 171 24 172 25
rect 172 24 173 25
rect 173 24 174 25
rect 174 24 175 25
rect 175 24 176 25
rect 176 24 177 25
rect 177 24 178 25
rect 194 24 195 25
rect 195 24 196 25
rect 196 24 197 25
rect 197 24 198 25
rect 198 24 199 25
rect 199 24 200 25
rect 200 24 201 25
rect 201 24 202 25
rect 217 24 218 25
rect 218 24 219 25
rect 219 24 220 25
rect 220 24 221 25
rect 264 24 265 25
rect 265 24 266 25
rect 266 24 267 25
rect 267 24 268 25
rect 268 24 269 25
rect 269 24 270 25
rect 270 24 271 25
rect 271 24 272 25
rect 272 24 273 25
rect 9 23 10 24
rect 10 23 11 24
rect 11 23 12 24
rect 12 23 13 24
rect 13 23 14 24
rect 14 23 15 24
rect 15 23 16 24
rect 34 23 35 24
rect 35 23 36 24
rect 36 23 37 24
rect 37 23 38 24
rect 38 23 39 24
rect 39 23 40 24
rect 40 23 41 24
rect 54 23 55 24
rect 55 23 56 24
rect 56 23 57 24
rect 57 23 58 24
rect 58 23 59 24
rect 59 23 60 24
rect 60 23 61 24
rect 72 23 73 24
rect 73 23 74 24
rect 74 23 75 24
rect 75 23 76 24
rect 76 23 77 24
rect 77 23 78 24
rect 78 23 79 24
rect 79 23 80 24
rect 91 23 92 24
rect 92 23 93 24
rect 93 23 94 24
rect 94 23 95 24
rect 125 23 126 24
rect 126 23 127 24
rect 127 23 128 24
rect 128 23 129 24
rect 129 23 130 24
rect 130 23 131 24
rect 131 23 132 24
rect 132 23 133 24
rect 133 23 134 24
rect 147 23 148 24
rect 148 23 149 24
rect 149 23 150 24
rect 150 23 151 24
rect 169 23 170 24
rect 170 23 171 24
rect 171 23 172 24
rect 172 23 173 24
rect 173 23 174 24
rect 174 23 175 24
rect 175 23 176 24
rect 176 23 177 24
rect 195 23 196 24
rect 196 23 197 24
rect 197 23 198 24
rect 198 23 199 24
rect 199 23 200 24
rect 200 23 201 24
rect 201 23 202 24
rect 202 23 203 24
rect 216 23 217 24
rect 217 23 218 24
rect 218 23 219 24
rect 219 23 220 24
rect 265 23 266 24
rect 266 23 267 24
rect 267 23 268 24
rect 268 23 269 24
rect 269 23 270 24
rect 270 23 271 24
rect 271 23 272 24
rect 9 22 10 23
rect 10 22 11 23
rect 11 22 12 23
rect 12 22 13 23
rect 13 22 14 23
rect 14 22 15 23
rect 15 22 16 23
rect 33 22 34 23
rect 34 22 35 23
rect 35 22 36 23
rect 36 22 37 23
rect 37 22 38 23
rect 38 22 39 23
rect 39 22 40 23
rect 40 22 41 23
rect 55 22 56 23
rect 56 22 57 23
rect 57 22 58 23
rect 58 22 59 23
rect 59 22 60 23
rect 60 22 61 23
rect 61 22 62 23
rect 71 22 72 23
rect 72 22 73 23
rect 73 22 74 23
rect 74 22 75 23
rect 75 22 76 23
rect 76 22 77 23
rect 77 22 78 23
rect 78 22 79 23
rect 79 22 80 23
rect 90 22 91 23
rect 91 22 92 23
rect 92 22 93 23
rect 93 22 94 23
rect 94 22 95 23
rect 125 22 126 23
rect 126 22 127 23
rect 127 22 128 23
rect 128 22 129 23
rect 129 22 130 23
rect 130 22 131 23
rect 131 22 132 23
rect 132 22 133 23
rect 133 22 134 23
rect 134 22 135 23
rect 146 22 147 23
rect 147 22 148 23
rect 148 22 149 23
rect 149 22 150 23
rect 170 22 171 23
rect 171 22 172 23
rect 172 22 173 23
rect 173 22 174 23
rect 174 22 175 23
rect 175 22 176 23
rect 176 22 177 23
rect 195 22 196 23
rect 196 22 197 23
rect 197 22 198 23
rect 198 22 199 23
rect 199 22 200 23
rect 200 22 201 23
rect 201 22 202 23
rect 202 22 203 23
rect 203 22 204 23
rect 204 22 205 23
rect 215 22 216 23
rect 216 22 217 23
rect 217 22 218 23
rect 218 22 219 23
rect 265 22 266 23
rect 266 22 267 23
rect 267 22 268 23
rect 268 22 269 23
rect 269 22 270 23
rect 270 22 271 23
rect 271 22 272 23
rect 9 21 10 22
rect 10 21 11 22
rect 11 21 12 22
rect 12 21 13 22
rect 13 21 14 22
rect 14 21 15 22
rect 15 21 16 22
rect 31 21 32 22
rect 32 21 33 22
rect 33 21 34 22
rect 34 21 35 22
rect 35 21 36 22
rect 36 21 37 22
rect 37 21 38 22
rect 38 21 39 22
rect 39 21 40 22
rect 55 21 56 22
rect 56 21 57 22
rect 57 21 58 22
rect 58 21 59 22
rect 59 21 60 22
rect 60 21 61 22
rect 61 21 62 22
rect 62 21 63 22
rect 71 21 72 22
rect 72 21 73 22
rect 73 21 74 22
rect 74 21 75 22
rect 75 21 76 22
rect 76 21 77 22
rect 77 21 78 22
rect 78 21 79 22
rect 79 21 80 22
rect 90 21 91 22
rect 91 21 92 22
rect 92 21 93 22
rect 93 21 94 22
rect 94 21 95 22
rect 95 21 96 22
rect 96 21 97 22
rect 97 21 98 22
rect 126 21 127 22
rect 127 21 128 22
rect 128 21 129 22
rect 129 21 130 22
rect 130 21 131 22
rect 131 21 132 22
rect 132 21 133 22
rect 133 21 134 22
rect 134 21 135 22
rect 135 21 136 22
rect 136 21 137 22
rect 143 21 144 22
rect 144 21 145 22
rect 145 21 146 22
rect 146 21 147 22
rect 147 21 148 22
rect 148 21 149 22
rect 170 21 171 22
rect 171 21 172 22
rect 172 21 173 22
rect 173 21 174 22
rect 174 21 175 22
rect 175 21 176 22
rect 176 21 177 22
rect 195 21 196 22
rect 196 21 197 22
rect 197 21 198 22
rect 198 21 199 22
rect 199 21 200 22
rect 200 21 201 22
rect 201 21 202 22
rect 202 21 203 22
rect 203 21 204 22
rect 204 21 205 22
rect 205 21 206 22
rect 213 21 214 22
rect 214 21 215 22
rect 215 21 216 22
rect 216 21 217 22
rect 217 21 218 22
rect 265 21 266 22
rect 266 21 267 22
rect 267 21 268 22
rect 268 21 269 22
rect 269 21 270 22
rect 270 21 271 22
rect 271 21 272 22
rect 9 20 10 21
rect 10 20 11 21
rect 11 20 12 21
rect 12 20 13 21
rect 13 20 14 21
rect 14 20 15 21
rect 15 20 16 21
rect 30 20 31 21
rect 31 20 32 21
rect 32 20 33 21
rect 33 20 34 21
rect 34 20 35 21
rect 35 20 36 21
rect 36 20 37 21
rect 37 20 38 21
rect 38 20 39 21
rect 55 20 56 21
rect 56 20 57 21
rect 57 20 58 21
rect 58 20 59 21
rect 59 20 60 21
rect 60 20 61 21
rect 61 20 62 21
rect 62 20 63 21
rect 63 20 64 21
rect 69 20 70 21
rect 70 20 71 21
rect 71 20 72 21
rect 73 20 74 21
rect 74 20 75 21
rect 75 20 76 21
rect 76 20 77 21
rect 77 20 78 21
rect 78 20 79 21
rect 79 20 80 21
rect 80 20 81 21
rect 90 20 91 21
rect 91 20 92 21
rect 92 20 93 21
rect 93 20 94 21
rect 94 20 95 21
rect 95 20 96 21
rect 96 20 97 21
rect 97 20 98 21
rect 98 20 99 21
rect 99 20 100 21
rect 100 20 101 21
rect 101 20 102 21
rect 102 20 103 21
rect 103 20 104 21
rect 104 20 105 21
rect 105 20 106 21
rect 106 20 107 21
rect 107 20 108 21
rect 108 20 109 21
rect 109 20 110 21
rect 110 20 111 21
rect 127 20 128 21
rect 128 20 129 21
rect 129 20 130 21
rect 130 20 131 21
rect 131 20 132 21
rect 132 20 133 21
rect 133 20 134 21
rect 134 20 135 21
rect 135 20 136 21
rect 136 20 137 21
rect 137 20 138 21
rect 138 20 139 21
rect 139 20 140 21
rect 140 20 141 21
rect 141 20 142 21
rect 142 20 143 21
rect 143 20 144 21
rect 144 20 145 21
rect 145 20 146 21
rect 146 20 147 21
rect 147 20 148 21
rect 148 20 149 21
rect 171 20 172 21
rect 172 20 173 21
rect 173 20 174 21
rect 174 20 175 21
rect 175 20 176 21
rect 196 20 197 21
rect 197 20 198 21
rect 198 20 199 21
rect 199 20 200 21
rect 200 20 201 21
rect 201 20 202 21
rect 202 20 203 21
rect 203 20 204 21
rect 204 20 205 21
rect 205 20 206 21
rect 206 20 207 21
rect 207 20 208 21
rect 208 20 209 21
rect 209 20 210 21
rect 210 20 211 21
rect 211 20 212 21
rect 212 20 213 21
rect 213 20 214 21
rect 214 20 215 21
rect 215 20 216 21
rect 216 20 217 21
rect 217 20 218 21
rect 266 20 267 21
rect 267 20 268 21
rect 268 20 269 21
rect 269 20 270 21
rect 270 20 271 21
rect 8 19 9 20
rect 9 19 10 20
rect 10 19 11 20
rect 11 19 12 20
rect 12 19 13 20
rect 13 19 14 20
rect 14 19 15 20
rect 15 19 16 20
rect 16 19 17 20
rect 17 19 18 20
rect 27 19 28 20
rect 28 19 29 20
rect 29 19 30 20
rect 30 19 31 20
rect 31 19 32 20
rect 32 19 33 20
rect 33 19 34 20
rect 34 19 35 20
rect 35 19 36 20
rect 36 19 37 20
rect 37 19 38 20
rect 55 19 56 20
rect 56 19 57 20
rect 57 19 58 20
rect 58 19 59 20
rect 59 19 60 20
rect 60 19 61 20
rect 61 19 62 20
rect 62 19 63 20
rect 63 19 64 20
rect 64 19 65 20
rect 65 19 66 20
rect 66 19 67 20
rect 67 19 68 20
rect 68 19 69 20
rect 69 19 70 20
rect 70 19 71 20
rect 71 19 72 20
rect 73 19 74 20
rect 74 19 75 20
rect 75 19 76 20
rect 76 19 77 20
rect 77 19 78 20
rect 78 19 79 20
rect 79 19 80 20
rect 80 19 81 20
rect 81 19 82 20
rect 82 19 83 20
rect 83 19 84 20
rect 90 19 91 20
rect 91 19 92 20
rect 92 19 93 20
rect 93 19 94 20
rect 94 19 95 20
rect 95 19 96 20
rect 96 19 97 20
rect 97 19 98 20
rect 98 19 99 20
rect 99 19 100 20
rect 100 19 101 20
rect 101 19 102 20
rect 102 19 103 20
rect 103 19 104 20
rect 104 19 105 20
rect 105 19 106 20
rect 106 19 107 20
rect 107 19 108 20
rect 108 19 109 20
rect 109 19 110 20
rect 110 19 111 20
rect 111 19 112 20
rect 112 19 113 20
rect 113 19 114 20
rect 114 19 115 20
rect 128 19 129 20
rect 129 19 130 20
rect 130 19 131 20
rect 131 19 132 20
rect 132 19 133 20
rect 133 19 134 20
rect 134 19 135 20
rect 135 19 136 20
rect 136 19 137 20
rect 137 19 138 20
rect 138 19 139 20
rect 139 19 140 20
rect 140 19 141 20
rect 141 19 142 20
rect 142 19 143 20
rect 143 19 144 20
rect 144 19 145 20
rect 145 19 146 20
rect 146 19 147 20
rect 147 19 148 20
rect 171 19 172 20
rect 172 19 173 20
rect 173 19 174 20
rect 174 19 175 20
rect 175 19 176 20
rect 197 19 198 20
rect 198 19 199 20
rect 199 19 200 20
rect 200 19 201 20
rect 201 19 202 20
rect 202 19 203 20
rect 203 19 204 20
rect 204 19 205 20
rect 205 19 206 20
rect 206 19 207 20
rect 207 19 208 20
rect 208 19 209 20
rect 209 19 210 20
rect 210 19 211 20
rect 211 19 212 20
rect 212 19 213 20
rect 213 19 214 20
rect 214 19 215 20
rect 215 19 216 20
rect 216 19 217 20
rect 266 19 267 20
rect 267 19 268 20
rect 268 19 269 20
rect 269 19 270 20
rect 270 19 271 20
rect 7 18 8 19
rect 8 18 9 19
rect 9 18 10 19
rect 10 18 11 19
rect 11 18 12 19
rect 12 18 13 19
rect 13 18 14 19
rect 14 18 15 19
rect 15 18 16 19
rect 16 18 17 19
rect 17 18 18 19
rect 18 18 19 19
rect 19 18 20 19
rect 20 18 21 19
rect 21 18 22 19
rect 22 18 23 19
rect 23 18 24 19
rect 24 18 25 19
rect 25 18 26 19
rect 26 18 27 19
rect 27 18 28 19
rect 28 18 29 19
rect 29 18 30 19
rect 30 18 31 19
rect 31 18 32 19
rect 32 18 33 19
rect 33 18 34 19
rect 34 18 35 19
rect 35 18 36 19
rect 36 18 37 19
rect 56 18 57 19
rect 57 18 58 19
rect 58 18 59 19
rect 59 18 60 19
rect 60 18 61 19
rect 61 18 62 19
rect 62 18 63 19
rect 63 18 64 19
rect 64 18 65 19
rect 65 18 66 19
rect 66 18 67 19
rect 67 18 68 19
rect 68 18 69 19
rect 69 18 70 19
rect 70 18 71 19
rect 73 18 74 19
rect 74 18 75 19
rect 75 18 76 19
rect 76 18 77 19
rect 77 18 78 19
rect 78 18 79 19
rect 79 18 80 19
rect 80 18 81 19
rect 81 18 82 19
rect 90 18 91 19
rect 91 18 92 19
rect 92 18 93 19
rect 93 18 94 19
rect 94 18 95 19
rect 95 18 96 19
rect 96 18 97 19
rect 97 18 98 19
rect 98 18 99 19
rect 99 18 100 19
rect 100 18 101 19
rect 101 18 102 19
rect 102 18 103 19
rect 103 18 104 19
rect 104 18 105 19
rect 105 18 106 19
rect 106 18 107 19
rect 107 18 108 19
rect 108 18 109 19
rect 109 18 110 19
rect 110 18 111 19
rect 111 18 112 19
rect 112 18 113 19
rect 113 18 114 19
rect 114 18 115 19
rect 115 18 116 19
rect 129 18 130 19
rect 130 18 131 19
rect 131 18 132 19
rect 132 18 133 19
rect 133 18 134 19
rect 134 18 135 19
rect 135 18 136 19
rect 136 18 137 19
rect 137 18 138 19
rect 138 18 139 19
rect 139 18 140 19
rect 140 18 141 19
rect 141 18 142 19
rect 142 18 143 19
rect 143 18 144 19
rect 144 18 145 19
rect 145 18 146 19
rect 171 18 172 19
rect 172 18 173 19
rect 173 18 174 19
rect 174 18 175 19
rect 175 18 176 19
rect 198 18 199 19
rect 199 18 200 19
rect 200 18 201 19
rect 201 18 202 19
rect 202 18 203 19
rect 203 18 204 19
rect 204 18 205 19
rect 205 18 206 19
rect 206 18 207 19
rect 207 18 208 19
rect 208 18 209 19
rect 209 18 210 19
rect 210 18 211 19
rect 211 18 212 19
rect 212 18 213 19
rect 213 18 214 19
rect 214 18 215 19
rect 266 18 267 19
rect 267 18 268 19
rect 268 18 269 19
rect 269 18 270 19
rect 1 17 2 18
rect 2 17 3 18
rect 3 17 4 18
rect 4 17 5 18
rect 5 17 6 18
rect 6 17 7 18
rect 7 17 8 18
rect 8 17 9 18
rect 9 17 10 18
rect 10 17 11 18
rect 11 17 12 18
rect 12 17 13 18
rect 13 17 14 18
rect 14 17 15 18
rect 15 17 16 18
rect 16 17 17 18
rect 17 17 18 18
rect 18 17 19 18
rect 19 17 20 18
rect 20 17 21 18
rect 21 17 22 18
rect 22 17 23 18
rect 23 17 24 18
rect 24 17 25 18
rect 25 17 26 18
rect 26 17 27 18
rect 27 17 28 18
rect 28 17 29 18
rect 29 17 30 18
rect 30 17 31 18
rect 31 17 32 18
rect 32 17 33 18
rect 33 17 34 18
rect 34 17 35 18
rect 57 17 58 18
rect 58 17 59 18
rect 59 17 60 18
rect 60 17 61 18
rect 61 17 62 18
rect 62 17 63 18
rect 63 17 64 18
rect 64 17 65 18
rect 65 17 66 18
rect 66 17 67 18
rect 67 17 68 18
rect 68 17 69 18
rect 69 17 70 18
rect 73 17 74 18
rect 74 17 75 18
rect 75 17 76 18
rect 76 17 77 18
rect 77 17 78 18
rect 78 17 79 18
rect 79 17 80 18
rect 92 17 93 18
rect 93 17 94 18
rect 94 17 95 18
rect 95 17 96 18
rect 96 17 97 18
rect 97 17 98 18
rect 98 17 99 18
rect 99 17 100 18
rect 100 17 101 18
rect 101 17 102 18
rect 102 17 103 18
rect 103 17 104 18
rect 104 17 105 18
rect 105 17 106 18
rect 106 17 107 18
rect 107 17 108 18
rect 108 17 109 18
rect 109 17 110 18
rect 110 17 111 18
rect 111 17 112 18
rect 112 17 113 18
rect 113 17 114 18
rect 114 17 115 18
rect 115 17 116 18
rect 116 17 117 18
rect 130 17 131 18
rect 131 17 132 18
rect 132 17 133 18
rect 133 17 134 18
rect 134 17 135 18
rect 135 17 136 18
rect 136 17 137 18
rect 137 17 138 18
rect 138 17 139 18
rect 139 17 140 18
rect 140 17 141 18
rect 141 17 142 18
rect 142 17 143 18
rect 143 17 144 18
rect 144 17 145 18
rect 172 17 173 18
rect 173 17 174 18
rect 174 17 175 18
rect 199 17 200 18
rect 200 17 201 18
rect 201 17 202 18
rect 202 17 203 18
rect 203 17 204 18
rect 204 17 205 18
rect 205 17 206 18
rect 206 17 207 18
rect 207 17 208 18
rect 208 17 209 18
rect 209 17 210 18
rect 210 17 211 18
rect 211 17 212 18
rect 212 17 213 18
rect 213 17 214 18
rect 267 17 268 18
rect 268 17 269 18
rect 269 17 270 18
rect 1 16 2 17
rect 3 16 4 17
rect 5 16 6 17
rect 6 16 7 17
rect 8 16 9 17
rect 10 16 11 17
rect 11 16 12 17
rect 13 16 14 17
rect 15 16 16 17
rect 16 16 17 17
rect 18 16 19 17
rect 20 16 21 17
rect 21 16 22 17
rect 23 16 24 17
rect 25 16 26 17
rect 26 16 27 17
rect 28 16 29 17
rect 30 16 31 17
rect 59 16 60 17
rect 60 16 61 17
rect 61 16 62 17
rect 62 16 63 17
rect 63 16 64 17
rect 64 16 65 17
rect 65 16 66 17
rect 67 16 68 17
rect 73 16 74 17
rect 74 16 75 17
rect 76 16 77 17
rect 93 16 94 17
rect 94 16 95 17
rect 95 16 96 17
rect 97 16 98 17
rect 98 16 99 17
rect 99 16 100 17
rect 100 16 101 17
rect 101 16 102 17
rect 102 16 103 17
rect 103 16 104 17
rect 104 16 105 17
rect 105 16 106 17
rect 106 16 107 17
rect 107 16 108 17
rect 108 16 109 17
rect 109 16 110 17
rect 110 16 111 17
rect 111 16 112 17
rect 112 16 113 17
rect 113 16 114 17
rect 114 16 115 17
rect 115 16 116 17
rect 116 16 117 17
rect 131 16 132 17
rect 133 16 134 17
rect 134 16 135 17
rect 135 16 136 17
rect 136 16 137 17
rect 137 16 138 17
rect 138 16 139 17
rect 139 16 140 17
rect 140 16 141 17
rect 142 16 143 17
rect 171 16 172 17
rect 172 16