magic
tech  scmos
timestamp 777777777
<< metal1 >>
rect 15 42 16 43
rect 28 42 29 43
rect 29 42 30 43
rect 30 42 31 43
rect 31 42 32 43
rect 32 42 33 43
rect 33 42 34 43
rect 34 42 35 43
rect 38 42 39 43
rect 39 42 40 43
rect 40 42 41 43
rect 41 42 42 43
rect 42 42 43 43
rect 43 42 44 43
rect 44 42 45 43
rect 45 42 46 43
rect 46 42 47 43
rect 47 42 48 43
rect 48 42 49 43
rect 58 42 59 43
rect 59 42 60 43
rect 60 42 61 43
rect 61 42 62 43
rect 62 42 63 43
rect 63 42 64 43
rect 64 42 65 43
rect 68 42 69 43
rect 69 42 70 43
rect 70 42 71 43
rect 71 42 72 43
rect 72 42 73 43
rect 73 42 74 43
rect 80 42 81 43
rect 81 42 82 43
rect 82 42 83 43
rect 83 42 84 43
rect 189 42 190 43
rect 190 42 191 43
rect 251 42 252 43
rect 252 42 253 43
rect 253 42 254 43
rect 15 41 16 42
rect 28 41 29 42
rect 29 41 30 42
rect 30 41 31 42
rect 31 41 32 42
rect 32 41 33 42
rect 33 41 34 42
rect 34 41 35 42
rect 38 41 39 42
rect 39 41 40 42
rect 40 41 41 42
rect 41 41 42 42
rect 42 41 43 42
rect 43 41 44 42
rect 44 41 45 42
rect 45 41 46 42
rect 46 41 47 42
rect 47 41 48 42
rect 48 41 49 42
rect 58 41 59 42
rect 59 41 60 42
rect 60 41 61 42
rect 61 41 62 42
rect 62 41 63 42
rect 63 41 64 42
rect 64 41 65 42
rect 68 41 69 42
rect 69 41 70 42
rect 70 41 71 42
rect 71 41 72 42
rect 72 41 73 42
rect 73 41 74 42
rect 80 41 81 42
rect 81 41 82 42
rect 82 41 83 42
rect 83 41 84 42
rect 189 41 190 42
rect 190 41 191 42
rect 251 41 252 42
rect 252 41 253 42
rect 253 41 254 42
rect 15 40 16 41
rect 16 40 17 41
rect 30 40 31 41
rect 31 40 32 41
rect 32 40 33 41
rect 33 40 34 41
rect 40 40 41 41
rect 44 40 45 41
rect 45 40 46 41
rect 46 40 47 41
rect 57 40 58 41
rect 58 40 59 41
rect 59 40 60 41
rect 62 40 63 41
rect 63 40 64 41
rect 64 40 65 41
rect 69 40 70 41
rect 70 40 71 41
rect 71 40 72 41
rect 72 40 73 41
rect 81 40 82 41
rect 82 40 83 41
rect 83 40 84 41
rect 184 40 185 41
rect 189 40 190 41
rect 190 40 191 41
rect 252 40 253 41
rect 253 40 254 41
rect 15 39 16 40
rect 16 39 17 40
rect 30 39 31 40
rect 31 39 32 40
rect 32 39 33 40
rect 33 39 34 40
rect 40 39 41 40
rect 44 39 45 40
rect 45 39 46 40
rect 46 39 47 40
rect 57 39 58 40
rect 58 39 59 40
rect 59 39 60 40
rect 62 39 63 40
rect 63 39 64 40
rect 64 39 65 40
rect 69 39 70 40
rect 70 39 71 40
rect 71 39 72 40
rect 72 39 73 40
rect 81 39 82 40
rect 82 39 83 40
rect 83 39 84 40
rect 184 39 185 40
rect 189 39 190 40
rect 190 39 191 40
rect 252 39 253 40
rect 253 39 254 40
rect 15 38 16 39
rect 16 38 17 39
rect 30 38 31 39
rect 31 38 32 39
rect 32 38 33 39
rect 33 38 34 39
rect 44 38 45 39
rect 45 38 46 39
rect 46 38 47 39
rect 56 38 57 39
rect 57 38 58 39
rect 58 38 59 39
rect 63 38 64 39
rect 64 38 65 39
rect 69 38 70 39
rect 70 38 71 39
rect 71 38 72 39
rect 72 38 73 39
rect 81 38 82 39
rect 82 38 83 39
rect 83 38 84 39
rect 183 38 184 39
rect 184 38 185 39
rect 189 38 190 39
rect 190 38 191 39
rect 252 38 253 39
rect 253 38 254 39
rect 15 37 16 38
rect 16 37 17 38
rect 30 37 31 38
rect 31 37 32 38
rect 32 37 33 38
rect 33 37 34 38
rect 44 37 45 38
rect 45 37 46 38
rect 46 37 47 38
rect 56 37 57 38
rect 57 37 58 38
rect 58 37 59 38
rect 63 37 64 38
rect 64 37 65 38
rect 69 37 70 38
rect 70 37 71 38
rect 71 37 72 38
rect 72 37 73 38
rect 81 37 82 38
rect 82 37 83 38
rect 83 37 84 38
rect 183 37 184 38
rect 184 37 185 38
rect 189 37 190 38
rect 190 37 191 38
rect 252 37 253 38
rect 253 37 254 38
rect 14 36 15 37
rect 15 36 16 37
rect 16 36 17 37
rect 31 36 32 37
rect 32 36 33 37
rect 33 36 34 37
rect 44 36 45 37
rect 45 36 46 37
rect 46 36 47 37
rect 56 36 57 37
rect 57 36 58 37
rect 58 36 59 37
rect 64 36 65 37
rect 69 36 70 37
rect 70 36 71 37
rect 71 36 72 37
rect 72 36 73 37
rect 81 36 82 37
rect 82 36 83 37
rect 83 36 84 37
rect 183 36 184 37
rect 184 36 185 37
rect 252 36 253 37
rect 253 36 254 37
rect 14 35 15 36
rect 15 35 16 36
rect 16 35 17 36
rect 31 35 32 36
rect 32 35 33 36
rect 33 35 34 36
rect 44 35 45 36
rect 45 35 46 36
rect 46 35 47 36
rect 56 35 57 36
rect 57 35 58 36
rect 58 35 59 36
rect 64 35 65 36
rect 69 35 70 36
rect 70 35 71 36
rect 71 35 72 36
rect 72 35 73 36
rect 81 35 82 36
rect 82 35 83 36
rect 83 35 84 36
rect 183 35 184 36
rect 184 35 185 36
rect 252 35 253 36
rect 253 35 254 36
rect 14 34 15 35
rect 15 34 16 35
rect 16 34 17 35
rect 31 34 32 35
rect 32 34 33 35
rect 33 34 34 35
rect 39 34 40 35
rect 44 34 45 35
rect 45 34 46 35
rect 46 34 47 35
rect 56 34 57 35
rect 57 34 58 35
rect 58 34 59 35
rect 59 34 60 35
rect 64 34 65 35
rect 69 34 70 35
rect 70 34 71 35
rect 71 34 72 35
rect 72 34 73 35
rect 81 34 82 35
rect 82 34 83 35
rect 83 34 84 35
rect 182 34 183 35
rect 183 34 184 35
rect 184 34 185 35
rect 252 34 253 35
rect 253 34 254 35
rect 14 33 15 34
rect 15 33 16 34
rect 16 33 17 34
rect 31 33 32 34
rect 32 33 33 34
rect 33 33 34 34
rect 39 33 40 34
rect 44 33 45 34
rect 45 33 46 34
rect 46 33 47 34
rect 56 33 57 34
rect 57 33 58 34
rect 58 33 59 34
rect 59 33 60 34
rect 64 33 65 34
rect 69 33 70 34
rect 70 33 71 34
rect 71 33 72 34
rect 72 33 73 34
rect 81 33 82 34
rect 82 33 83 34
rect 83 33 84 34
rect 182 33 183 34
rect 183 33 184 34
rect 184 33 185 34
rect 252 33 253 34
rect 253 33 254 34
rect 13 32 14 33
rect 15 32 16 33
rect 16 32 17 33
rect 17 32 18 33
rect 31 32 32 33
rect 32 32 33 33
rect 33 32 34 33
rect 39 32 40 33
rect 44 32 45 33
rect 45 32 46 33
rect 46 32 47 33
rect 56 32 57 33
rect 57 32 58 33
rect 58 32 59 33
rect 59 32 60 33
rect 60 32 61 33
rect 69 32 70 33
rect 70 32 71 33
rect 71 32 72 33
rect 72 32 73 33
rect 81 32 82 33
rect 82 32 83 33
rect 83 32 84 33
rect 89 32 90 33
rect 90 32 91 33
rect 91 32 92 33
rect 98 32 99 33
rect 99 32 100 33
rect 100 32 101 33
rect 101 32 102 33
rect 102 32 103 33
rect 103 32 104 33
rect 104 32 105 33
rect 109 32 110 33
rect 110 32 111 33
rect 111 32 112 33
rect 124 32 125 33
rect 125 32 126 33
rect 126 32 127 33
rect 127 32 128 33
rect 128 32 129 33
rect 129 32 130 33
rect 135 32 136 33
rect 136 32 137 33
rect 137 32 138 33
rect 141 32 142 33
rect 142 32 143 33
rect 143 32 144 33
rect 144 32 145 33
rect 146 32 147 33
rect 147 32 148 33
rect 148 32 149 33
rect 149 32 150 33
rect 155 32 156 33
rect 156 32 157 33
rect 157 32 158 33
rect 162 32 163 33
rect 163 32 164 33
rect 164 32 165 33
rect 166 32 167 33
rect 167 32 168 33
rect 168 32 169 33
rect 173 32 174 33
rect 174 32 175 33
rect 175 32 176 33
rect 176 32 177 33
rect 181 32 182 33
rect 182 32 183 33
rect 183 32 184 33
rect 184 32 185 33
rect 185 32 186 33
rect 186 32 187 33
rect 188 32 189 33
rect 189 32 190 33
rect 190 32 191 33
rect 196 32 197 33
rect 197 32 198 33
rect 198 32 199 33
rect 199 32 200 33
rect 204 32 205 33
rect 205 32 206 33
rect 206 32 207 33
rect 207 32 208 33
rect 208 32 209 33
rect 209 32 210 33
rect 210 32 211 33
rect 211 32 212 33
rect 212 32 213 33
rect 220 32 221 33
rect 221 32 222 33
rect 222 32 223 33
rect 223 32 224 33
rect 224 32 225 33
rect 225 32 226 33
rect 226 32 227 33
rect 227 32 228 33
rect 233 32 234 33
rect 234 32 235 33
rect 235 32 236 33
rect 236 32 237 33
rect 244 32 245 33
rect 245 32 246 33
rect 246 32 247 33
rect 247 32 248 33
rect 252 32 253 33
rect 253 32 254 33
rect 256 32 257 33
rect 257 32 258 33
rect 258 32 259 33
rect 259 32 260 33
rect 264 32 265 33
rect 265 32 266 33
rect 266 32 267 33
rect 267 32 268 33
rect 274 32 275 33
rect 275 32 276 33
rect 276 32 277 33
rect 277 32 278 33
rect 278 32 279 33
rect 279 32 280 33
rect 285 32 286 33
rect 286 32 287 33
rect 287 32 288 33
rect 13 31 14 32
rect 16 31 17 32
rect 17 31 18 32
rect 32 31 33 32
rect 33 31 34 32
rect 34 31 35 32
rect 38 31 39 32
rect 44 31 45 32
rect 45 31 46 32
rect 46 31 47 32
rect 56 31 57 32
rect 57 31 58 32
rect 58 31 59 32
rect 59 31 60 32
rect 60 31 61 32
rect 61 31 62 32
rect 69 31 70 32
rect 70 31 71 32
rect 71 31 72 32
rect 72 31 73 32
rect 81 31 82 32
rect 82 31 83 32
rect 83 31 84 32
rect 87 31 88 32
rect 88 31 89 32
rect 89 31 90 32
rect 91 31 92 32
rect 92 31 93 32
rect 93 31 94 32
rect 97 31 98 32
rect 98 31 99 32
rect 99 31 100 32
rect 101 31 102 32
rect 102 31 103 32
rect 107 31 108 32
rect 108 31 109 32
rect 109 31 110 32
rect 112 31 113 32
rect 113 31 114 32
rect 123 31 124 32
rect 124 31 125 32
rect 126 31 127 32
rect 127 31 128 32
rect 128 31 129 32
rect 133 31 134 32
rect 134 31 135 32
rect 137 31 138 32
rect 138 31 139 32
rect 142 31 143 32
rect 143 31 144 32
rect 144 31 145 32
rect 145 31 146 32
rect 148 31 149 32
rect 149 31 150 32
rect 150 31 151 32
rect 153 31 154 32
rect 154 31 155 32
rect 157 31 158 32
rect 158 31 159 32
rect 163 31 164 32
rect 164 31 165 32
rect 165 31 166 32
rect 166 31 167 32
rect 167 31 168 32
rect 168 31 169 32
rect 172 31 173 32
rect 173 31 174 32
rect 176 31 177 32
rect 177 31 178 32
rect 178 31 179 32
rect 182 31 183 32
rect 183 31 184 32
rect 184 31 185 32
rect 189 31 190 32
rect 190 31 191 32
rect 195 31 196 32
rect 196 31 197 32
rect 199 31 200 32
rect 200 31 201 32
rect 201 31 202 32
rect 205 31 206 32
rect 206 31 207 32
rect 207 31 208 32
rect 211 31 212 32
rect 212 31 213 32
rect 221 31 222 32
rect 222 31 223 32
rect 223 31 224 32
rect 226 31 227 32
rect 227 31 228 32
rect 228 31 229 32
rect 232 31 233 32
rect 233 31 234 32
rect 236 31 237 32
rect 237 31 238 32
rect 238 31 239 32
rect 243 31 244 32
rect 244 31 245 32
rect 247 31 248 32
rect 248 31 249 32
rect 252 31 253 32
rect 253 31 254 32
rect 257 31 258 32
rect 263 31 264 32
rect 267 31 268 32
rect 268 31 269 32
rect 273 31 274 32
rect 274 31 275 32
rect 276 31 277 32
rect 277 31 278 32
rect 278 31 279 32
rect 283 31 284 32
rect 284 31 285 32
rect 287 31 288 32
rect 288 31 289 32
rect 13 30 14 31
rect 16 30 17 31
rect 17 30 18 31
rect 32 30 33 31
rect 33 30 34 31
rect 34 30 35 31
rect 38 30 39 31
rect 44 30 45 31
rect 45 30 46 31
rect 46 30 47 31
rect 56 30 57 31
rect 57 30 58 31
rect 58 30 59 31
rect 59 30 60 31
rect 60 30 61 31
rect 61 30 62 31
rect 69 30 70 31
rect 70 30 71 31
rect 71 30 72 31
rect 72 30 73 31
rect 81 30 82 31
rect 82 30 83 31
rect 83 30 84 31
rect 87 30 88 31
rect 88 30 89 31
rect 89 30 90 31
rect 91 30 92 31
rect 92 30 93 31
rect 93 30 94 31
rect 97 30 98 31
rect 98 30 99 31
rect 99 30 100 31
rect 101 30 102 31
rect 102 30 103 31
rect 107 30 108 31
rect 108 30 109 31
rect 109 30 110 31
rect 112 30 113 31
rect 113 30 114 31
rect 123 30 124 31
rect 124 30 125 31
rect 126 30 127 31
rect 127 30 128 31
rect 128 30 129 31
rect 133 30 134 31
rect 134 30 135 31
rect 137 30 138 31
rect 138 30 139 31
rect 142 30 143 31
rect 143 30 144 31
rect 144 30 145 31
rect 145 30 146 31
rect 148 30 149 31
rect 149 30 150 31
rect 150 30 151 31
rect 153 30 154 31
rect 154 30 155 31
rect 157 30 158 31
rect 158 30 159 31
rect 163 30 164 31
rect 164 30 165 31
rect 165 30 166 31
rect 166 30 167 31
rect 167 30 168 31
rect 168 30 169 31
rect 172 30 173 31
rect 173 30 174 31
rect 176 30 177 31
rect 177 30 178 31
rect 178 30 179 31
rect 182 30 183 31
rect 183 30 184 31
rect 184 30 185 31
rect 189 30 190 31
rect 190 30 191 31
rect 195 30 196 31
rect 196 30 197 31
rect 199 30 200 31
rect 200 30 201 31
rect 201 30 202 31
rect 205 30 206 31
rect 206 30 207 31
rect 207 30 208 31
rect 211 30 212 31
rect 212 30 213 31
rect 221 30 222 31
rect 222 30 223 31
rect 223 30 224 31
rect 226 30 227 31
rect 227 30 228 31
rect 228 30 229 31
rect 232 30 233 31
rect 233 30 234 31
rect 236 30 237 31
rect 237 30 238 31
rect 238 30 239 31
rect 243 30 244 31
rect 244 30 245 31
rect 247 30 248 31
rect 248 30 249 31
rect 252 30 253 31
rect 253 30 254 31
rect 257 30 258 31
rect 263 30 264 31
rect 267 30 268 31
rect 268 30 269 31
rect 273 30 274 31
rect 274 30 275 31
rect 276 30 277 31
rect 277 30 278 31
rect 278 30 279 31
rect 283 30 284 31
rect 284 30 285 31
rect 287 30 288 31
rect 288 30 289 31
rect 12 29 13 30
rect 16 29 17 30
rect 17 29 18 30
rect 32 29 33 30
rect 33 29 34 30
rect 34 29 35 30
rect 38 29 39 30
rect 44 29 45 30
rect 45 29 46 30
rect 46 29 47 30
rect 57 29 58 30
rect 58 29 59 30
rect 59 29 60 30
rect 60 29 61 30
rect 61 29 62 30
rect 62 29 63 30
rect 63 29 64 30
rect 69 29 70 30
rect 70 29 71 30
rect 71 29 72 30
rect 72 29 73 30
rect 81 29 82 30
rect 82 29 83 30
rect 83 29 84 30
rect 87 29 88 30
rect 88 29 89 30
rect 92 29 93 30
rect 93 29 94 30
rect 96 29 97 30
rect 97 29 98 30
rect 98 29 99 30
rect 101 29 102 30
rect 102 29 103 30
rect 103 29 104 30
rect 107 29 108 30
rect 108 29 109 30
rect 112 29 113 30
rect 113 29 114 30
rect 122 29 123 30
rect 123 29 124 30
rect 127 29 128 30
rect 128 29 129 30
rect 133 29 134 30
rect 134 29 135 30
rect 137 29 138 30
rect 138 29 139 30
rect 139 29 140 30
rect 142 29 143 30
rect 143 29 144 30
rect 144 29 145 30
rect 148 29 149 30
rect 149 29 150 30
rect 150 29 151 30
rect 153 29 154 30
rect 154 29 155 30
rect 157 29 158 30
rect 158 29 159 30
rect 159 29 160 30
rect 163 29 164 30
rect 164 29 165 30
rect 165 29 166 30
rect 167 29 168 30
rect 168 29 169 30
rect 171 29 172 30
rect 172 29 173 30
rect 173 29 174 30
rect 176 29 177 30
rect 177 29 178 30
rect 178 29 179 30
rect 182 29 183 30
rect 183 29 184 30
rect 184 29 185 30
rect 189 29 190 30
rect 190 29 191 30
rect 195 29 196 30
rect 200 29 201 30
rect 201 29 202 30
rect 205 29 206 30
rect 206 29 207 30
rect 207 29 208 30
rect 211 29 212 30
rect 212 29 213 30
rect 221 29 222 30
rect 222 29 223 30
rect 223 29 224 30
rect 227 29 228 30
rect 228 29 229 30
rect 231 29 232 30
rect 232 29 233 30
rect 233 29 234 30
rect 236 29 237 30
rect 237 29 238 30
rect 238 29 239 30
rect 242 29 243 30
rect 243 29 244 30
rect 247 29 248 30
rect 248 29 249 30
rect 252 29 253 30
rect 253 29 254 30
rect 256 29 257 30
rect 257 29 258 30
rect 262 29 263 30
rect 263 29 264 30
rect 267 29 268 30
rect 268 29 269 30
rect 272 29 273 30
rect 273 29 274 30
rect 274 29 275 30
rect 277 29 278 30
rect 278 29 279 30
rect 279 29 280 30
rect 283 29 284 30
rect 284 29 285 30
rect 287 29 288 30
rect 288 29 289 30
rect 289 29 290 30
rect 12 28 13 29
rect 16 28 17 29
rect 17 28 18 29
rect 32 28 33 29
rect 33 28 34 29
rect 34 28 35 29
rect 38 28 39 29
rect 44 28 45 29
rect 45 28 46 29
rect 46 28 47 29
rect 57 28 58 29
rect 58 28 59 29
rect 59 28 60 29
rect 60 28 61 29
rect 61 28 62 29
rect 62 28 63 29
rect 63 28 64 29
rect 69 28 70 29
rect 70 28 71 29
rect 71 28 72 29
rect 72 28 73 29
rect 81 28 82 29
rect 82 28 83 29
rect 83 28 84 29
rect 87 28 88 29
rect 88 28 89 29
rect 92 28 93 29
rect 93 28 94 29
rect 96 28 97 29
rect 97 28 98 29
rect 98 28 99 29
rect 101 28 102 29
rect 102 28 103 29
rect 103 28 104 29
rect 107 28 108 29
rect 108 28 109 29
rect 112 28 113 29
rect 113 28 114 29
rect 122 28 123 29
rect 123 28 124 29
rect 127 28 128 29
rect 128 28 129 29
rect 133 28 134 29
rect 134 28 135 29
rect 137 28 138 29
rect 138 28 139 29
rect 139 28 140 29
rect 142 28 143 29
rect 143 28 144 29
rect 144 28 145 29
rect 148 28 149 29
rect 149 28 150 29
rect 150 28 151 29
rect 153 28 154 29
rect 154 28 155 29
rect 157 28 158 29
rect 158 28 159 29
rect 159 28 160 29
rect 163 28 164 29
rect 164 28 165 29
rect 165 28 166 29
rect 167 28 168 29
rect 168 28 169 29
rect 171 28 172 29
rect 172 28 173 29
rect 173 28 174 29
rect 176 28 177 29
rect 177 28 178 29
rect 178 28 179 29
rect 182 28 183 29
rect 183 28 184 29
rect 184 28 185 29
rect 189 28 190 29
rect 190 28 191 29
rect 195 28 196 29
rect 200 28 201 29
rect 201 28 202 29
rect 205 28 206 29
rect 206 28 207 29
rect 207 28 208 29
rect 211 28 212 29
rect 212 28 213 29
rect 221 28 222 29
rect 222 28 223 29
rect 223 28 224 29
rect 227 28 228 29
rect 228 28 229 29
rect 231 28 232 29
rect 232 28 233 29
rect 233 28 234 29
rect 236 28 237 29
rect 237 28 238 29
rect 238 28 239 29
rect 242 28 243 29
rect 243 28 244 29
rect 247 28 248 29
rect 248 28 249 29
rect 252 28 253 29
rect 253 28 254 29
rect 256 28 257 29
rect 257 28 258 29
rect 262 28 263 29
rect 263 28 264 29
rect 267 28 268 29
rect 268 28 269 29
rect 272 28 273 29
rect 273 28 274 29
rect 274 28 275 29
rect 277 28 278 29
rect 278 28 279 29
rect 279 28 280 29
rect 283 28 284 29
rect 284 28 285 29
rect 287 28 288 29
rect 288 28 289 29
rect 289 28 290 29
rect 12 27 13 28
rect 17 27 18 28
rect 18 27 19 28
rect 33 27 34 28
rect 34 27 35 28
rect 35 27 36 28
rect 37 27 38 28
rect 44 27 45 28
rect 45 27 46 28
rect 46 27 47 28
rect 58 27 59 28
rect 59 27 60 28
rect 60 27 61 28
rect 61 27 62 28
rect 62 27 63 28
rect 63 27 64 28
rect 64 27 65 28
rect 69 27 70 28
rect 70 27 71 28
rect 71 27 72 28
rect 72 27 73 28
rect 81 27 82 28
rect 82 27 83 28
rect 83 27 84 28
rect 86 27 87 28
rect 87 27 88 28
rect 88 27 89 28
rect 92 27 93 28
rect 93 27 94 28
rect 94 27 95 28
rect 96 27 97 28
rect 97 27 98 28
rect 98 27 99 28
rect 101 27 102 28
rect 102 27 103 28
rect 103 27 104 28
rect 107 27 108 28
rect 108 27 109 28
rect 112 27 113 28
rect 113 27 114 28
rect 114 27 115 28
rect 122 27 123 28
rect 123 27 124 28
rect 127 27 128 28
rect 128 27 129 28
rect 132 27 133 28
rect 133 27 134 28
rect 134 27 135 28
rect 137 27 138 28
rect 138 27 139 28
rect 139 27 140 28
rect 142 27 143 28
rect 143 27 144 28
rect 144 27 145 28
rect 148 27 149 28
rect 149 27 150 28
rect 150 27 151 28
rect 152 27 153 28
rect 153 27 154 28
rect 154 27 155 28
rect 157 27 158 28
rect 158 27 159 28
rect 159 27 160 28
rect 163 27 164 28
rect 164 27 165 28
rect 171 27 172 28
rect 172 27 173 28
rect 173 27 174 28
rect 176 27 177 28
rect 177 27 178 28
rect 178 27 179 28
rect 182 27 183 28
rect 183 27 184 28
rect 184 27 185 28
rect 189 27 190 28
rect 190 27 191 28
rect 194 27 195 28
rect 195 27 196 28
rect 200 27 201 28
rect 201 27 202 28
rect 205 27 206 28
rect 206 27 207 28
rect 207 27 208 28
rect 211 27 212 28
rect 212 27 213 28
rect 221 27 222 28
rect 222 27 223 28
rect 223 27 224 28
rect 227 27 228 28
rect 228 27 229 28
rect 229 27 230 28
rect 231 27 232 28
rect 232 27 233 28
rect 233 27 234 28
rect 236 27 237 28
rect 237 27 238 28
rect 238 27 239 28
rect 241 27 242 28
rect 242 27 243 28
rect 243 27 244 28
rect 247 27 248 28
rect 248 27 249 28
rect 252 27 253 28
rect 253 27 254 28
rect 256 27 257 28
rect 262 27 263 28
rect 263 27 264 28
rect 267 27 268 28
rect 268 27 269 28
rect 272 27 273 28
rect 273 27 274 28
rect 274 27 275 28
rect 277 27 278 28
rect 278 27 279 28
rect 279 27 280 28
rect 282 27 283 28
rect 283 27 284 28
rect 284 27 285 28
rect 287 27 288 28
rect 288 27 289 28
rect 289 27 290 28
rect 12 26 13 27
rect 17 26 18 27
rect 18 26 19 27
rect 33 26 34 27
rect 34 26 35 27
rect 35 26 36 27
rect 37 26 38 27
rect 44 26 45 27
rect 45 26 46 27
rect 46 26 47 27
rect 58 26 59 27
rect 59 26 60 27
rect 60 26 61 27
rect 61 26 62 27
rect 62 26 63 27
rect 63 26 64 27
rect 64 26 65 27
rect 69 26 70 27
rect 70 26 71 27
rect 71 26 72 27
rect 72 26 73 27
rect 81 26 82 27
rect 82 26 83 27
rect 83 26 84 27
rect 86 26 87 27
rect 87 26 88 27
rect 88 26 89 27
rect 92 26 93 27
rect 93 26 94 27
rect 94 26 95 27
rect 96 26 97 27
rect 97 26 98 27
rect 98 26 99 27
rect 101 26 102 27
rect 102 26 103 27
rect 103 26 104 27
rect 107 26 108 27
rect 108 26 109 27
rect 112 26 113 27
rect 113 26 114 27
rect 114 26 115 27
rect 122 26 123 27
rect 123 26 124 27
rect 127 26 128 27
rect 128 26 129 27
rect 132 26 133 27
rect 133 26 134 27
rect 134 26 135 27
rect 137 26 138 27
rect 138 26 139 27
rect 139 26 140 27
rect 142 26 143 27
rect 143 26 144 27
rect 144 26 145 27
rect 148 26 149 27
rect 149 26 150 27
rect 150 26 151 27
rect 152 26 153 27
rect 153 26 154 27
rect 154 26 155 27
rect 157 26 158 27
rect 158 26 159 27
rect 159 26 160 27
rect 163 26 164 27
rect 164 26 165 27
rect 171 26 172 27
rect 172 26 173 27
rect 173 26 174 27
rect 176 26 177 27
rect 177 26 178 27
rect 178 26 179 27
rect 182 26 183 27
rect 183 26 184 27
rect 184 26 185 27
rect 189 26 190 27
rect 190 26 191 27
rect 194 26 195 27
rect 195 26 196 27
rect 200 26 201 27
rect 201 26 202 27
rect 205 26 206 27
rect 206 26 207 27
rect 207 26 208 27
rect 211 26 212 27
rect 212 26 213 27
rect 221 26 222 27
rect 222 26 223 27
rect 223 26 224 27
rect 227 26 228 27
rect 228 26 229 27
rect 229 26 230 27
rect 231 26 232 27
rect 232 26 233 27
rect 233 26 234 27
rect 236 26 237 27
rect 237 26 238 27
rect 238 26 239 27
rect 241 26 242 27
rect 242 26 243 27
rect 243 26 244 27
rect 247 26 248 27
rect 248 26 249 27
rect 252 26 253 27
rect 253 26 254 27
rect 256 26 257 27
rect 262 26 263 27
rect 263 26 264 27
rect 267 26 268 27
rect 268 26 269 27
rect 272 26 273 27
rect 273 26 274 27
rect 274 26 275 27
rect 277 26 278 27
rect 278 26 279 27
rect 279 26 280 27
rect 282 26 283 27
rect 283 26 284 27
rect 284 26 285 27
rect 287 26 288 27
rect 288 26 289 27
rect 289 26 290 27
rect 12 25 13 26
rect 17 25 18 26
rect 18 25 19 26
rect 33 25 34 26
rect 34 25 35 26
rect 35 25 36 26
rect 37 25 38 26
rect 44 25 45 26
rect 45 25 46 26
rect 46 25 47 26
rect 60 25 61 26
rect 61 25 62 26
rect 62 25 63 26
rect 63 25 64 26
rect 64 25 65 26
rect 65 25 66 26
rect 69 25 70 26
rect 70 25 71 26
rect 71 25 72 26
rect 72 25 73 26
rect 81 25 82 26
rect 82 25 83 26
rect 83 25 84 26
rect 86 25 87 26
rect 87 25 88 26
rect 88 25 89 26
rect 92 25 93 26
rect 93 25 94 26
rect 94 25 95 26
rect 96 25 97 26
rect 97 25 98 26
rect 98 25 99 26
rect 101 25 102 26
rect 102 25 103 26
rect 103 25 104 26
rect 107 25 108 26
rect 108 25 109 26
rect 112 25 113 26
rect 113 25 114 26
rect 114 25 115 26
rect 122 25 123 26
rect 123 25 124 26
rect 127 25 128 26
rect 128 25 129 26
rect 132 25 133 26
rect 133 25 134 26
rect 134 25 135 26
rect 135 25 136 26
rect 136 25 137 26
rect 137 25 138 26
rect 138 25 139 26
rect 139 25 140 26
rect 142 25 143 26
rect 143 25 144 26
rect 144 25 145 26
rect 148 25 149 26
rect 149 25 150 26
rect 150 25 151 26
rect 152 25 153 26
rect 153 25 154 26
rect 154 25 155 26
rect 155 25 156 26
rect 156 25 157 26
rect 157 25 158 26
rect 158 25 159 26
rect 159 25 160 26
rect 163 25 164 26
rect 164 25 165 26
rect 171 25 172 26
rect 172 25 173 26
rect 173 25 174 26
rect 176 25 177 26
rect 177 25 178 26
rect 178 25 179 26
rect 182 25 183 26
rect 183 25 184 26
rect 184 25 185 26
rect 189 25 190 26
rect 190 25 191 26
rect 194 25 195 26
rect 195 25 196 26
rect 200 25 201 26
rect 201 25 202 26
rect 205 25 206 26
rect 206 25 207 26
rect 207 25 208 26
rect 211 25 212 26
rect 212 25 213 26
rect 221 25 222 26
rect 222 25 223 26
rect 223 25 224 26
rect 227 25 228 26
rect 228 25 229 26
rect 229 25 230 26
rect 231 25 232 26
rect 232 25 233 26
rect 233 25 234 26
rect 236 25 237 26
rect 237 25 238 26
rect 238 25 239 26
rect 241 25 242 26
rect 242 25 243 26
rect 243 25 244 26
rect 252 25 253 26
rect 253 25 254 26
rect 255 25 256 26
rect 256 25 257 26
rect 262 25 263 26
rect 263 25 264 26
rect 267 25 268 26
rect 268 25 269 26
rect 272 25 273 26
rect 273 25 274 26
rect 274 25 275 26
rect 277 25 278 26
rect 278 25 279 26
rect 279 25 280 26
rect 282 25 283 26
rect 283 25 284 26
rect 284 25 285 26
rect 285 25 286 26
rect 286 25 287 26
rect 287 25 288 26
rect 288 25 289 26
rect 289 25 290 26
rect 12 24 13 25
rect 17 24 18 25
rect 18 24 19 25
rect 33 24 34 25
rect 34 24 35 25
rect 35 24 36 25
rect 37 24 38 25
rect 44 24 45 25
rect 45 24 46 25
rect 46 24 47 25
rect 60 24 61 25
rect 61 24 62 25
rect 62 24 63 25
rect 63 24 64 25
rect 64 24 65 25
rect 65 24 66 25
rect 69 24 70 25
rect 70 24 71 25
rect 71 24 72 25
rect 72 24 73 25
rect 81 24 82 25
rect 82 24 83 25
rect 83 24 84 25
rect 86 24 87 25
rect 87 24 88 25
rect 88 24 89 25
rect 92 24 93 25
rect 93 24 94 25
rect 94 24 95 25
rect 96 24 97 25
rect 97 24 98 25
rect 98 24 99 25
rect 101 24 102 25
rect 102 24 103 25
rect 103 24 104 25
rect 107 24 108 25
rect 108 24 109 25
rect 112 24 113 25
rect 113 24 114 25
rect 114 24 115 25
rect 122 24 123 25
rect 123 24 124 25
rect 127 24 128 25
rect 128 24 129 25
rect 132 24 133 25
rect 133 24 134 25
rect 134 24 135 25
rect 135 24 136 25
rect 136 24 137 25
rect 137 24 138 25
rect 138 24 139 25
rect 139 24 140 25
rect 142 24 143 25
rect 143 24 144 25
rect 144 24 145 25
rect 148 24 149 25
rect 149 24 150 25
rect 150 24 151 25
rect 152 24 153 25
rect 153 24 154 25
rect 154 24 155 25
rect 155 24 156 25
rect 156 24 157 25
rect 157 24 158 25
rect 158 24 159 25
rect 159 24 160 25
rect 163 24 164 25
rect 164 24 165 25
rect 171 24 172 25
rect 172 24 173 25
rect 173 24 174 25
rect 176 24 177 25
rect 177 24 178 25
rect 178 24 179 25
rect 182 24 183 25
rect 183 24 184 25
rect 184 24 185 25
rect 189 24 190 25
rect 190 24 191 25
rect 194 24 195 25
rect 195 24 196 25
rect 200 24 201 25
rect 201 24 202 25
rect 205 24 206 25
rect 206 24 207 25
rect 207 24 208 25
rect 211 24 212 25
rect 212 24 213 25
rect 221 24 222 25
rect 222 24 223 25
rect 223 24 224 25
rect 227 24 228 25
rect 228 24 229 25
rect 229 24 230 25
rect 231 24 232 25
rect 232 24 233 25
rect 233 24 234 25
rect 236 24 237 25
rect 237 24 238 25
rect 238 24 239 25
rect 241 24 242 25
rect 242 24 243 25
rect 243 24 244 25
rect 252 24 253 25
rect 253 24 254 25
rect 255 24 256 25
rect 256 24 257 25
rect 262 24 263 25
rect 263 24 264 25
rect 267 24 268 25
rect 268 24 269 25
rect 272 24 273 25
rect 273 24 274 25
rect 274 24 275 25
rect 277 24 278 25
rect 278 24 279 25
rect 279 24 280 25
rect 282 24 283 25
rect 283 24 284 25
rect 284 24 285 25
rect 285 24 286 25
rect 286 24 287 25
rect 287 24 288 25
rect 288 24 289 25
rect 289 24 290 25
rect 12 23 13 24
rect 13 23 14 24
rect 14 23 15 24
rect 15 23 16 24
rect 16 23 17 24
rect 17 23 18 24
rect 18 23 19 24
rect 19 23 20 24
rect 34 23 35 24
rect 35 23 36 24
rect 36 23 37 24
rect 37 23 38 24
rect 44 23 45 24
rect 45 23 46 24
rect 46 23 47 24
rect 54 23 55 24
rect 56 23 57 24
rect 62 23 63 24
rect 63 23 64 24
rect 64 23 65 24
rect 65 23 66 24
rect 69 23 70 24
rect 70 23 71 24
rect 71 23 72 24
rect 72 23 73 24
rect 81 23 82 24
rect 82 23 83 24
rect 83 23 84 24
rect 86 23 87 24
rect 87 23 88 24
rect 88 23 89 24
rect 92 23 93 24
rect 93 23 94 24
rect 94 23 95 24
rect 96 23 97 24
rect 97 23 98 24
rect 98 23 99 24
rect 101 23 102 24
rect 102 23 103 24
rect 103 23 104 24
rect 107 23 108 24
rect 108 23 109 24
rect 112 23 113 24
rect 113 23 114 24
rect 114 23 115 24
rect 122 23 123 24
rect 123 23 124 24
rect 127 23 128 24
rect 128 23 129 24
rect 132 23 133 24
rect 133 23 134 24
rect 134 23 135 24
rect 142 23 143 24
rect 143 23 144 24
rect 144 23 145 24
rect 148 23 149 24
rect 149 23 150 24
rect 150 23 151 24
rect 152 23 153 24
rect 153 23 154 24
rect 154 23 155 24
rect 163 23 164 24
rect 164 23 165 24
rect 174 23 175 24
rect 175 23 176 24
rect 176 23 177 24
rect 177 23 178 24
rect 178 23 179 24
rect 182 23 183 24
rect 183 23 184 24
rect 184 23 185 24
rect 189 23 190 24
rect 190 23 191 24
rect 194 23 195 24
rect 195 23 196 24
rect 200 23 201 24
rect 201 23 202 24
rect 205 23 206 24
rect 206 23 207 24
rect 207 23 208 24
rect 211 23 212 24
rect 212 23 213 24
rect 221 23 222 24
rect 222 23 223 24
rect 223 23 224 24
rect 227 23 228 24
rect 228 23 229 24
rect 229 23 230 24
rect 234 23 235 24
rect 235 23 236 24
rect 236 23 237 24
rect 237 23 238 24
rect 238 23 239 24
rect 241 23 242 24
rect 242 23 243 24
rect 243 23 244 24
rect 252 23 253 24
rect 253 23 254 24
rect 254 23 255 24
rect 255 23 256 24
rect 256 23 257 24
rect 257 23 258 24
rect 264 23 265 24
rect 265 23 266 24
rect 266 23 267 24
rect 267 23 268 24
rect 268 23 269 24
rect 272 23 273 24
rect 273 23 274 24
rect 274 23 275 24
rect 277 23 278 24
rect 278 23 279 24
rect 279 23 280 24
rect 282 23 283 24
rect 283 23 284 24
rect 284 23 285 24
rect 12 22 13 23
rect 13 22 14 23
rect 14 22 15 23
rect 15 22 16 23
rect 16 22 17 23
rect 17 22 18 23
rect 18 22 19 23
rect 19 22 20 23
rect 34 22 35 23
rect 35 22 36 23
rect 36 22 37 23
rect 37 22 38 23
rect 44 22 45 23
rect 45 22 46 23
rect 46 22 47 23
rect 54 22 55 23
rect 56 22 57 23
rect 62 22 63 23
rect 63 22 64 23
rect 64 22 65 23
rect 65 22 66 23
rect 69 22 70 23
rect 70 22 71 23
rect 71 22 72 23
rect 72 22 73 23
rect 81 22 82 23
rect 82 22 83 23
rect 83 22 84 23
rect 86 22 87 23
rect 87 22 88 23
rect 88 22 89 23
rect 92 22 93 23
rect 93 22 94 23
rect 94 22 95 23
rect 96 22 97 23
rect 97 22 98 23
rect 98 22 99 23
rect 101 22 102 23
rect 102 22 103 23
rect 103 22 104 23
rect 107 22 108 23
rect 108 22 109 23
rect 112 22 113 23
rect 113 22 114 23
rect 114 22 115 23
rect 122 22 123 23
rect 123 22 124 23
rect 127 22 128 23
rect 128 22 129 23
rect 132 22 133 23
rect 133 22 134 23
rect 134 22 135 23
rect 142 22 143 23
rect 143 22 144 23
rect 144 22 145 23
rect 148 22 149 23
rect 149 22 150 23
rect 150 22 151 23
rect 152 22 153 23
rect 153 22 154 23
rect 154 22 155 23
rect 163 22 164 23
rect 164 22 165 23
rect 174 22 175 23
rect 175 22 176 23
rect 176 22 177 23
rect 177 22 178 23
rect 178 22 179 23
rect 182 22 183 23
rect 183 22 184 23
rect 184 22 185 23
rect 189 22 190 23
rect 190 22 191 23
rect 194 22 195 23
rect 195 22 196 23
rect 200 22 201 23
rect 201 22 202 23
rect 205 22 206 23
rect 206 22 207 23
rect 207 22 208 23
rect 211 22 212 23
rect 212 22 213 23
rect 221 22 222 23
rect 222 22 223 23
rect 223 22 224 23
rect 227 22 228 23
rect 228 22 229 23
rect 229 22 230 23
rect 234 22 235 23
rect 235 22 236 23
rect 236 22 237 23
rect 237 22 238 23
rect 238 22 239 23
rect 241 22 242 23
rect 242 22 243 23
rect 243 22 244 23
rect 252 22 253 23
rect 253 22 254 23
rect 254 22 255 23
rect 255 22 256 23
rect 256 22 257 23
rect 257 22 258 23
rect 264 22 265 23
rect 265 22 266 23
rect 266 22 267 23
rect 267 22 268 23
rect 268 22 269 23
rect 272 22 273 23
rect 273 22 274 23
rect 274 22 275 23
rect 277 22 278 23
rect 278 22 279 23
rect 279 22 280 23
rect 282 22 283 23
rect 283 22 284 23
rect 284 22 285 23
rect 17 21 18 22
rect 18 21 19 22
rect 19 21 20 22
rect 34 21 35 22
rect 35 21 36 22
rect 36 21 37 22
rect 44 21 45 22
rect 45 21 46 22
rect 46 21 47 22
rect 54 21 55 22
rect 56 21 57 22
rect 63 21 64 22
rect 64 21 65 22
rect 65 21 66 22
rect 69 21 70 22
rect 70 21 71 22
rect 71 21 72 22
rect 72 21 73 22
rect 81 21 82 22
rect 82 21 83 22
rect 83 21 84 22
rect 86 21 87 22
rect 87 21 88 22
rect 88 21 89 22
rect 92 21 93 22
rect 93 21 94 22
rect 94 21 95 22
rect 97 21 98 22
rect 98 21 99 22
rect 99 21 100 22
rect 101 21 102 22
rect 102 21 103 22
rect 107 21 108 22
rect 108 21 109 22
rect 112 21 113 22
rect 113 21 114 22
rect 114 21 115 22
rect 123 21 124 22
rect 124 21 125 22
rect 126 21 127 22
rect 127 21 128 22
rect 128 21 129 22
rect 132 21 133 22
rect 133 21 134 22
rect 134 21 135 22
rect 142 21 143 22
rect 143 21 144 22
rect 144 21 145 22
rect 148 21 149 22
rect 149 21 150 22
rect 150 21 151 22
rect 152 21 153 22
rect 153 21 154 22
rect 154 21 155 22
rect 163 21 164 22
rect 164 21 165 22
rect 172 21 173 22
rect 173 21 174 22
rect 176 21 177 22
rect 177 21 178 22
rect 178 21 179 22
rect 182 21 183 22
rect 183 21 184 22
rect 184 21 185 22
rect 189 21 190 22
rect 190 21 191 22
rect 194 21 195 22
rect 195 21 196 22
rect 200 21 201 22
rect 201 21 202 22
rect 205 21 206 22
rect 206 21 207 22
rect 207 21 208 22
rect 211 21 212 22
rect 212 21 213 22
rect 221 21 222 22
rect 222 21 223 22
rect 223 21 224 22
rect 227 21 228 22
rect 228 21 229 22
rect 229 21 230 22
rect 232 21 233 22
rect 233 21 234 22
rect 234 21 235 22
rect 236 21 237 22
rect 237 21 238 22
rect 238 21 239 22
rect 241 21 242 22
rect 242 21 243 22
rect 243 21 244 22
rect 252 21 253 22
rect 253 21 254 22
rect 255 21 256 22
rect 256 21 257 22
rect 257 21 258 22
rect 263 21 264 22
rect 264 21 265 22
rect 267 21 268 22
rect 268 21 269 22
rect 273 21 274 22
rect 274 21 275 22
rect 276 21 277 22
rect 277 21 278 22
rect 278 21 279 22
rect 282 21 283 22
rect 283 21 284 22
rect 284 21 285 22
rect 17 20 18 21
rect 18 20 19 21
rect 19 20 20 21
rect 34 20 35 21
rect 35 20 36 21
rect 36 20 37 21
rect 44 20 45 21
rect 45 20 46 21
rect 46 20 47 21
rect 54 20 55 21
rect 56 20 57 21
rect 63 20 64 21
rect 64 20 65 21
rect 65 20 66 21
rect 69 20 70 21
rect 70 20 71 21
rect 71 20 72 21
rect 72 20 73 21
rect 81 20 82 21
rect 82 20 83 21
rect 83 20 84 21
rect 86 20 87 21
rect 87 20 88 21
rect 88 20 89 21
rect 92 20 93 21
rect 93 20 94 21
rect 94 20 95 21
rect 97 20 98 21
rect 98 20 99 21
rect 99 20 100 21
rect 101 20 102 21
rect 102 20 103 21
rect 107 20 108 21
rect 108 20 109 21
rect 112 20 113 21
rect 113 20 114 21
rect 114 20 115 21
rect 123 20 124 21
rect 124 20 125 21
rect 126 20 127 21
rect 127 20 128 21
rect 128 20 129 21
rect 132 20 133 21
rect 133 20 134 21
rect 134 20 135 21
rect 142 20 143 21
rect 143 20 144 21
rect 144 20 145 21
rect 148 20 149 21
rect 149 20 150 21
rect 150 20 151 21
rect 152 20 153 21
rect 153 20 154 21
rect 154 20 155 21
rect 163 20 164 21
rect 164 20 165 21
rect 172 20 173 21
rect 173 20 174 21
rect 176 20 177 21
rect 177 20 178 21
rect 178 20 179 21
rect 182 20 183 21
rect 183 20 184 21
rect 184 20 185 21
rect 189 20 190 21
rect 190 20 191 21
rect 194 20 195 21
rect 195 20 196 21
rect 200 20 201 21
rect 201 20 202 21
rect 205 20 206 21
rect 206 20 207 21
rect 207 20 208 21
rect 211 20 212 21
rect 212 20 213 21
rect 221 20 222 21
rect 222 20 223 21
rect 223 20 224 21
rect 227 20 228 21
rect 228 20 229 21
rect 229 20 230 21
rect 232 20 233 21
rect 233 20 234 21
rect 234 20 235 21
rect 236 20 237 21
rect 237 20 238 21
rect 238 20 239 21
rect 241 20 242 21
rect 242 20 243 21
rect 243 20 244 21
rect 252 20 253 21
rect 253 20 254 21
rect 255 20 256 21
rect 256 20 257 21
rect 257 20 258 21
rect 263 20 264 21
rect 264 20 265 21
rect 267 20 268 21
rect 268 20 269 21
rect 273 20 274 21
rect 274 20 275 21
rect 276 20 277 21
rect 277 20 278 21
rect 278 20 279 21
rect 282 20 283 21
rect 283 20 284 21
rect 284 20 285 21
rect 11 19 12 20
rect 17 19 18 20
rect 18 19 19 20
rect 19 19 20 20
rect 20 19 21 20
rect 34 19 35 20
rect 35 19 36 20
rect 36 19 37 20
rect 44 19 45 20
rect 45 19 46 20
rect 46 19 47 20
rect 53 19 54 20
rect 54 19 55 20
rect 56 19 57 20
rect 63 19 64 20
rect 64 19 65 20
rect 65 19 66 20
rect 69 19 70 20
rect 70 19 71 20
rect 71 19 72 20
rect 72 19 73 20
rect 81 19 82 20
rect 82 19 83 20
rect 83 19 84 20
rect 86 19 87 20
rect 87 19 88 20
rect 88 19 89 20
rect 92 19 93 20
rect 93 19 94 20
rect 94 19 95 20
rect 99 19 100 20
rect 100 19 101 20
rect 101 19 102 20
rect 107 19 108 20
rect 108 19 109 20
rect 112 19 113 20
rect 113 19 114 20
rect 114 19 115 20
rect 124 19 125 20
rect 125 19 126 20
rect 126 19 127 20
rect 127 19 128 20
rect 132 19 133 20
rect 133 19 134 20
rect 134 19 135 20
rect 142 19 143 20
rect 143 19 144 20
rect 144 19 145 20
rect 148 19 149 20
rect 149 19 150 20
rect 150 19 151 20
rect 152 19 153 20
rect 153 19 154 20
rect 154 19 155 20
rect 163 19 164 20
rect 164 19 165 20
rect 171 19 172 20
rect 172 19 173 20
rect 173 19 174 20
rect 176 19 177 20
rect 177 19 178 20
rect 178 19 179 20
rect 182 19 183 20
rect 183 19 184 20
rect 184 19 185 20
rect 189 19 190 20
rect 190 19 191 20
rect 194 19 195 20
rect 195 19 196 20
rect 200 19 201 20
rect 201 19 202 20
rect 205 19 206 20
rect 206 19 207 20
rect 207 19 208 20
rect 211 19 212 20
rect 212 19 213 20
rect 221 19 222 20
rect 222 19 223 20
rect 223 19 224 20
rect 227 19 228 20
rect 228 19 229 20
rect 229 19 230 20
rect 231 19 232 20
rect 232 19 233 20
rect 233 19 234 20
rect 236 19 237 20
rect 237 19 238 20
rect 238 19 239 20
rect 241 19 242 20
rect 242 19 243 20
rect 243 19 244 20
rect 244 19 245 20
rect 252 19 253 20
rect 253 19 254 20
rect 255 19 256 20
rect 256 19 257 20
rect 257 19 258 20
rect 262 19 263 20
rect 263 19 264 20
rect 267 19 268 20
rect 268 19 269 20
rect 275 19 276 20
rect 276 19 277 20
rect 277 19 278 20
rect 282 19 283 20
rect 283 19 284 20
rect 284 19 285 20
rect 11 18 12 19
rect 17 18 18 19
rect 18 18 19 19
rect 19 18 20 19
rect 20 18 21 19
rect 34 18 35 19
rect 35 18 36 19
rect 36 18 37 19
rect 44 18 45 19
rect 45 18 46 19
rect 46 18 47 19
rect 53 18 54 19
rect 54 18 55 19
rect 56 18 57 19
rect 63 18 64 19
rect 64 18 65 19
rect 65 18 66 19
rect 69 18 70 19
rect 70 18 71 19
rect 71 18 72 19
rect 72 18 73 19
rect 81 18 82 19
rect 82 18 83 19
rect 83 18 84 19
rect 86 18 87 19
rect 87 18 88 19
rect 88 18 89 19
rect 92 18 93 19
rect 93 18 94 19
rect 94 18 95 19
rect 99 18 100 19
rect 100 18 101 19
rect 101 18 102 19
rect 107 18 108 19
rect 108 18 109 19
rect 112 18 113 19
rect 113 18 114 19
rect 114 18 115 19
rect 124 18 125 19
rect 125 18 126 19
rect 126 18 127 19
rect 127 18 128 19
rect 132 18 133 19
rect 133 18 134 19
rect 134 18 135 19
rect 142 18 143 19
rect 143 18 144 19
rect 144 18 145 19
rect 148 18 149 19
rect 149 18 150 19
rect 150 18 151 19
rect 152 18 153 19
rect 153 18 154 19
rect 154 18 155 19
rect 163 18 164 19
rect 164 18 165 19
rect 171 18 172 19
rect 172 18 173 19
rect 173 18 174 19
rect 176 18 177 19
rect 177 18 178 19
rect 178 18 179 19
rect 182 18 183 19
rect 183 18 184 19
rect 184 18 185 19
rect 189 18 190 19
rect 190 18 191 19
rect 194 18 195 19
rect 195 18 196 19
rect 200 18 201 19
rect 201 18 202 19
rect 205 18 206 19
rect 206 18 207 19
rect 207 18 208 19
rect 211 18 212 19
rect 212 18 213 19
rect 221 18 222 19
rect 222 18 223 19
rect 223 18 224 19
rect 227 18 228 19
rect 228 18 229 19
rect 229 18 230 19
rect 231 18 232 19
rect 232 18 233 19
rect 233 18 234 19
rect 236 18 237 19
rect 237 18 238 19
rect 238 18 239 19
rect 241 18 242 19
rect 242 18 243 19
rect 243 18 244 19
rect 244 18 245 19
rect 252 18 253 19
rect 253 18 254 19
rect 255 18 256 19
rect 256 18 257 19
rect 257 18 258 19
rect 262 18 263 19
rect 263 18 264 19
rect 267 18 268 19
rect 268 18 269 19
rect 275 18 276 19
rect 276 18 277 19
rect 277 18 278 19
rect 282 18 283 19
rect 283 18 284 19
rect 284 18 285 19
rect 11 17 12 18
rect 17 17 18 18
rect 18 17 19 18
rect 19 17 20 18
rect 20 17 21 18
rect 34 17 35 18
rect 35 17 36 18
rect 44 17 45 18
rect 45 17 46 18
rect 46 17 47 18
rect 52 17 53 18
rect 53 17 54 18
rect 56 17 57 18
rect 57 17 58 18
rect 63 17 64 18
rect 64 17 65 18
rect 69 17 70 18
rect 70 17 71 18
rect 71 17 72 18
rect 72 17 73 18
rect 81 17 82 18
rect 82 17 83 18
rect 83 17 84 18
rect 87 17 88 18
rect 88 17 89 18
rect 92 17 93 18
rect 93 17 94 18
rect 97 17 98 18
rect 98 17 99 18
rect 107 17 108 18
rect 108 17 109 18
rect 112 17 113 18
rect 113 17 114 18
rect 123 17 124 18
rect 133 17 134 18
rect 134 17 135 18
rect 139 17 140 18
rect 142 17 143 18
rect 143 17 144 18
rect 144 17 145 18
rect 148 17 149 18
rect 149 17 150 18
rect 150 17 151 18
rect 153 17 154 18
rect 154 17 155 18
rect 155 17 156 18
rect 159 17 160 18
rect 163 17 164 18
rect 164 17 165 18
rect 171 17 172 18
rect 172 17 173 18
rect 173 17 174 18
rect 176 17 177 18
rect 177 17 178 18
rect 178 17 179 18
rect 182 17 183 18
rect 183 17 184 18
rect 184 17 185 18
rect 189 17 190 18
rect 190 17 191 18
rect 195 17 196 18
rect 200 17 201 18
rect 201 17 202 18
rect 205 17 206 18
rect 206 17 207 18
rect 207 17 208 18
rect 211 17 212 18
rect 212 17 213 18
rect 221 17 222 18
rect 222 17 223 18
rect 223 17 224 18
rect 227 17 228 18
rect 228 17 229 18
rect 231 17 232 18
rect 232 17 233 18
rect 233 17 234 18
rect 236 17 237 18
rect 237 17 238 18
rect 238 17 239 18
rect 242 17 243 18
rect 243 17 244 18
rect 244 17 245 18
rect 245 17 246 18
rect 248 17 249 18
rect 252 17 253 18
rect 253 17 254 18
rect 256 17 257 18
rect 257 17 258 18
rect 258 17 259 18
rect 262 17 263 18
rect 263 17 264 18
rect 267 17 268 18
rect 268 17 269 18
rect 273 17 274 18
rect 274 17 275 18
rect 283 17 284 18
rect 284 17 285 18
rect 285 17 286 18
rect 289 17 290 18
rect 11 16 12 17
rect 17 16 18 17
rect 18 16 19 17
rect 19 16 20 17
rect 20 16 21 17
rect 34 16 35 17
rect 35 16 36 17
rect 44 16 45 17
rect 45 16 46 17
rect 46 16 47 17
rect 52 16 53 17
rect 53 16 54 17
rect 56 16 57 17
rect 57 16 58 17
rect 63 16 64 17
rect 64 16 65 17
rect 69 16 70 17
rect 70 16 71 17
rect 71 16 72 17
rect 72 16 73 17
rect 81 16 82 17
rect 82 16 83 17
rect 83 16 84 17
rect 87 16 88 17
rect 88 16 89 17
rect 92 16 93 17
rect 93 16 94 17
rect 97 16 98 17
rect 98 16 99 17
rect 107 16 108 17
rect 108 16 109 17
rect 112 16 113 17
rect 113 16 114 17
rect 123 16 124 17
rect 133 16 134 17
rect 134 16 135 17
rect 139 16 140 17
rect 142 16 143 17
rect 143 16 144 17
rect 144 16 145 17
rect 148 16 149 17
rect 149 16 150 17
rect 150 16 151 17
rect 153 16 154 17
rect 154 16 155 17
rect 155 16 156 17
rect 159 16 160 17
rect 163 16 164 17
rect 164 16 165 17
rect 171 16 172 17
rect 172 16 173 17
rect 173 16 174 17
rect 176 16 177 17
rect 177 16 178 17
rect 178 16 179 17
rect 182 16 183 17
rect 183 16 184 17
rect 184 16 185 17
rect 189 16 190 17
rect 190 16 191 17
rect 195 16 196 17
rect 200 16 201 17
rect 201 16 202 17
rect 205 16 206 17
rect 206 16 207 17
rect 207 16 208 17
rect 211 16 212 17
rect 212 16 213 17
rect 221 16 222 17
rect 222 16 223 17
rect 223 16 224 17
rect 227 16 228 17
rect 228 16 229 17
rect 231 16 232 17
rect 232 16 233 17
rect 233 16 234 17
rect 236 16 237 17
rect 237 16 238 17
rect 238 16 239 17
rect 242 16 243 17
rect 243 16 244 17
rect 244 16 245 17
rect 245 16 246 17
rect 248 16 249 17
rect 252 16 253 17
rect 253 16 254 17
rect 256 16 257 17
rect 257 16 258 17
rect 258 16 259 17
rect 262 16 263 17
rect 263 16 264 17
rect 267 16 268 17
rect 268 16 269 17
rect 273 16 274 17
rect 274 16 275 17
rect 283 16 284 17
rect 284 16 285 17
rect 285 16 286 17
rect 289 16 290 17
rect 10 15 11 16
rect 11 15 12 16
rect 17 15 18 16
rect 18 15 19 16
rect 19 15 20 16
rect 20 15 21 16
rect 21 15 22 16
rect 34 15 35 16
rect 35 15 36 16
rect 44 15 45 16
rect 45 15 46 16
rect 46 15 47 16
rect 51 15 52 16
rect 52 15 53 16
rect 53 15 54 16
rect 56 15 57 16
rect 57 15 58 16
rect 58 15 59 16
rect 62 15 63 16
rect 63 15 64 16
rect 64 15 65 16
rect 69 15 70 16
rect 70 15 71 16
rect 71 15 72 16
rect 72 15 73 16
rect 81 15 82 16
rect 82 15 83 16
rect 83 15 84 16
rect 87 15 88 16
rect 88 15 89 16
rect 89 15 90 16
rect 91 15 92 16
rect 92 15 93 16
rect 93 15 94 16
rect 96 15 97 16
rect 97 15 98 16
rect 98 15 99 16
rect 107 15 108 16
rect 108 15 109 16
rect 109 15 110 16
rect 112 15 113 16
rect 113 15 114 16
rect 122 15 123 16
rect 123 15 124 16
rect 133 15 134 16
rect 134 15 135 16
rect 135 15 136 16
rect 136 15 137 16
rect 137 15 138 16
rect 138 15 139 16
rect 142 15 143 16
rect 143 15 144 16
rect 144 15 145 16
rect 148 15 149 16
rect 149 15 150 16
rect 150 15 151 16
rect 153 15 154 16
rect 154 15 155 16
rect 155 15 156 16
rect 156 15 157 16
rect 157 15 158 16
rect 158 15 159 16
rect 163 15 164 16
rect 164 15 165 16
rect 171 15 172 16
rect 172 15 173 16
rect 173 15 174 16
rect 174 15 175 16
rect 175 15 176 16
rect 176 15 177 16
rect 177 15 178 16
rect 178 15 179 16
rect 179 15 180 16
rect 182 15 183 16
rect 183 15 184 16
rect 184 15 185 16
rect 186 15 187 16
rect 189 15 190 16
rect 190 15 191 16
rect 195 15 196 16
rect 196 15 197 16
rect 199 15 200 16
rect 200 15 201 16
rect 201 15 202 16
rect 205 15 206 16
rect 206 15 207 16
rect 207 15 208 16
rect 211 15 212 16
rect 212 15 213 16
rect 221 15 222 16
rect 222 15 223 16
rect 223 15 224 16
rect 226 15 227 16
rect 227 15 228 16
rect 228 15 229 16
rect 231 15 232 16
rect 232 15 233 16
rect 233 15 234 16
rect 234 15 235 16
rect 235 15 236 16
rect 236 15 237 16
rect 237 15 238 16
rect 238 15 239 16
rect 239 15 240 16
rect 242 15 243 16
rect 243 15 244 16
rect 244 15 245 16
rect 245 15 246 16
rect 246 15 247 16
rect 247 15 248 16
rect 252 15 253 16
rect 253 15 254 16
rect 257 15 258 16
rect 258 15 259 16
rect 259 15 260 16
rect 262 15 263 16
rect 263 15 264 16
rect 264 15 265 16
rect 265 15 266 16
rect 266 15 267 16
rect 267 15 268 16
rect 268 15 269 16
rect 269 15 270 16
rect 272 15 273 16
rect 273 15 274 16
rect 274 15 275 16
rect 283 15 284 16
rect 284 15 285 16
rect 285 15 286 16
rect 286 15 287 16
rect 287 15 288 16
rect 288 15 289 16
rect 10 14 11 15
rect 11 14 12 15
rect 17 14 18 15
rect 18 14 19 15
rect 19 14 20 15
rect 20 14 21 15
rect 21 14 22 15
rect 34 14 35 15
rect 35 14 36 15
rect 44 14 45 15
rect 45 14 46 15
rect 46 14 47 15
rect 51 14 52 15
rect 52 14 53 15
rect 53 14 54 15
rect 56 14 57 15
rect 57 14 58 15
rect 58 14 59 15
rect 62 14 63 15
rect 63 14 64 15
rect 64 14 65 15
rect 69 14 70 15
rect 70 14 71 15
rect 71 14 72 15
rect 72 14 73 15
rect 81 14 82 15
rect 82 14 83 15
rect 83 14 84 15
rect 87 14 88 15
rect 88 14 89 15
rect 89 14 90 15
rect 91 14 92 15
rect 92 14 93 15
rect 93 14 94 15
rect 96 14 97 15
rect 97 14 98 15
rect 98 14 99 15
rect 107 14 108 15
rect 108 14 109 15
rect 109 14 110 15
rect 112 14 113 15
rect 113 14 114 15
rect 122 14 123 15
rect 123 14 124 15
rect 133 14 134 15
rect 134 14 135 15
rect 135 14 136 15
rect 136 14 137 15
rect 137 14 138 15
rect 138 14 139 15
rect 142 14 143 15
rect 143 14 144 15
rect 144 14 145 15
rect 148 14 149 15
rect 149 14 150 15
rect 150 14 151 15
rect 153 14 154 15
rect 154 14 155 15
rect 155 14 156 15
rect 156 14 157 15
rect 157 14 158 15
rect 158 14 159 15
rect 163 14 164 15
rect 164 14 165 15
rect 171 14 172 15
rect 172 14 173 15
rect 173 14 174 15
rect 174 14 175 15
rect 175 14 176 15
rect 176 14 177 15
rect 177 14 178 15
rect 178 14 179 15
rect 179 14 180 15
rect 182 14 183 15
rect 183 14 184 15
rect 184 14 185 15
rect 186 14 187 15
rect 189 14 190 15
rect 190 14 191 15
rect 195 14 196 15
rect 196 14 197 15
rect 199 14 200 15
rect 200 14 201 15
rect 201 14 202 15
rect 205 14 206 15
rect 206 14 207 15
rect 207 14 208 15
rect 211 14 212 15
rect 212 14 213 15
rect 221 14 222 15
rect 222 14 223 15
rect 223 14 224 15
rect 226 14 227 15
rect 227 14 228 15
rect 228 14 229 15
rect 231 14 232 15
rect 232 14 233 15
rect 233 14 234 15
rect 234 14 235 15
rect 235 14 236 15
rect 236 14 237 15
rect 237 14 238 15
rect 238 14 239 15
rect 239 14 240 15
rect 242 14 243 15
rect 243 14 244 15
rect 244 14 245 15
rect 245 14 246 15
rect 246 14 247 15
rect 247 14 248 15
rect 252 14 253 15
rect 253 14 254 15
rect 257 14 258 15
rect 258 14 259 15
rect 259 14 260 15
rect 262 14 263 15
rect 263 14 264 15
rect 264 14 265 15
rect 265 14 266 15
rect 266 14 267 15
rect 267 14 268 15
rect 268 14 269 15
rect 269 14 270 15
rect 272 14 273 15
rect 273 14 274 15
rect 274 14 275 15
rect 283 14 284 15
rect 284 14 285 15
rect 285 14 286 15
rect 286 14 287 15
rect 287 14 288 15
rect 288 14 289 15
rect 9 13 10 14
rect 10 13 11 14
rect 11 13 12 14
rect 12 13 13 14
rect 16 13 17 14
rect 17 13 18 14
rect 18 13 19 14
rect 19 13 20 14
rect 20 13 21 14
rect 21 13 22 14
rect 22 13 23 14
rect 34 13 35 14
rect 42 13 43 14
rect 43 13 44 14
rect 44 13 45 14
rect 45 13 46 14
rect 46 13 47 14
rect 47 13 48 14
rect 48 13 49 14
rect 49 13 50 14
rect 50 13 51 14
rect 51 13 52 14
rect 52 13 53 14
rect 53 13 54 14
rect 56 13 57 14
rect 59 13 60 14
rect 60 13 61 14
rect 61 13 62 14
rect 62 13 63 14
rect 68 13 69 14
rect 69 13 70 14
rect 70 13 71 14
rect 71 13 72 14
rect 72 13 73 14
rect 73 13 74 14
rect 80 13 81 14
rect 81 13 82 14
rect 82 13 83 14
rect 83 13 84 14
rect 89 13 90 14
rect 90 13 91 14
rect 91 13 92 14
rect 96 13 97 14
rect 97 13 98 14
rect 98 13 99 14
rect 99 13 100 14
rect 100 13 101 14
rect 101 13 102 14
rect 102 13 103 14
rect 103 13 104 14
rect 109 13 110 14
rect 110 13 111 14
rect 111 13 112 14
rect 122 13 123 14
rect 123 13 124 14
rect 124 13 125 14
rect 125 13 126 14
rect 126 13 127 14
rect 127 13 128 14
rect 128 13 129 14
rect 135 13 136 14
rect 136 13 137 14
rect 137 13 138 14
rect 141 13 142 14
rect 142 13 143 14
rect 143 13 144 14
rect 144 13 145 14
rect 145 13 146 14
rect 147 13 148 14
rect 148 13 149 14
rect 149 13 150 14
rect 150 13 151 14
rect 151 13 152 14
rect 155 13 156 14
rect 156 13 157 14
rect 157 13 158 14
rect 162 13 163 14
rect 163 13 164 14
rect 164 13 165 14
rect 165 13 166 14
rect 172 13 173 14
rect 173 13 174 14
rect 176 13 177 14
rect 177 13 178 14
rect 178 13 179 14
rect 183 13 184 14
rect 184 13 185 14
rect 185 13 186 14
rect 188 13 189 14
rect 189 13 190 14
rect 190 13 191 14
rect 191 13 192 14
rect 196 13 197 14
rect 197 13 198 14
rect 198 13 199 14
rect 199 13 200 14
rect 204 13 205 14
rect 205 13 206 14
rect 206 13 207 14
rect 207 13 208 14
rect 210 13 211 14
rect 211 13 212 14
rect 212 13 213 14
rect 213 13 214 14
rect 221 13 222 14
rect 222 13 223 14
rect 223 13 224 14
rect 224 13 225 14
rect 225 13 226 14
rect 226 13 227 14
rect 227 13 228 14
rect 232 13 233 14
rect 233 13 234 14
rect 234 13 235 14
rect 236 13 237 14
rect 237 13 238 14
rect 238 13 239 14
rect 244 13 245 14
rect 245 13 246 14
rect 246 13 247 14
rect 251 13 252 14
rect 252 13 253 14
rect 253 13 254 14
rect 254 13 255 14
rect 256 13 257 14
rect 257 13 258 14
rect 258 13 259 14
rect 259 13 260 14
rect 260 13 261 14
rect 263 13 264 14
rect 264 13 265 14
rect 267 13 268 14
rect 268 13 269 14
rect 272 13 273 14
rect 273 13 274 14
rect 274 13 275 14
rect 275 13 276 14
rect 276 13 277 14
rect 277 13 278 14
rect 278 13 279 14
rect 279 13 280 14
rect 285 13 286 14
rect 286 13 287 14
rect 287 13 288 14
rect 9 12 10 13
rect 10 12 11 13
rect 11 12 12 13
rect 12 12 13 13
rect 16 12 17 13
rect 17 12 18 13
rect 18 12 19 13
rect 19 12 20 13
rect 20 12 21 13
rect 21 12 22 13
rect 22 12 23 13
rect 34 12 35 13
rect 42 12 43 13
rect 43 12 44 13
rect 44 12 45 13
rect 45 12 46 13
rect 46 12 47 13
rect 47 12 48 13
rect 48 12 49 13
rect 49 12 50 13
rect 50 12 51 13
rect 51 12 52 13
rect 52 12 53 13
rect 53 12 54 13
rect 56 12 57 13
rect 59 12 60 13
rect 60 12 61 13
rect 61 12 62 13
rect 62 12 63 13
rect 68 12 69 13
rect 69 12 70 13
rect 70 12 71 13
rect 71 12 72 13
rect 72 12 73 13
rect 73 12 74 13
rect 80 12 81 13
rect 81 12 82 13
rect 82 12 83 13
rect 83 12 84 13
rect 89 12 90 13
rect 90 12 91 13
rect 91 12 92 13
rect 96 12 97 13
rect 97 12 98 13
rect 98 12 99 13
rect 99 12 100 13
rect 100 12 101 13
rect 101 12 102 13
rect 102 12 103 13
rect 103 12 104 13
rect 109 12 110 13
rect 110 12 111 13
rect 111 12 112 13
rect 122 12 123 13
rect 123 12 124 13
rect 124 12 125 13
rect 125 12 126 13
rect 126 12 127 13
rect 127 12 128 13
rect 128 12 129 13
rect 135 12 136 13
rect 136 12 137 13
rect 137 12 138 13
rect 141 12 142 13
rect 142 12 143 13
rect 143 12 144 13
rect 144 12 145 13
rect 145 12 146 13
rect 147 12 148 13
rect 148 12 149 13
rect 149 12 150 13
rect 150 12 151 13
rect 151 12 152 13
rect 155 12 156 13
rect 156 12 157 13
rect 157 12 158 13
rect 162 12 163 13
rect 163 12 164 13
rect 164 12 165 13
rect 165 12 166 13
rect 172 12 173 13
rect 173 12 174 13
rect 176 12 177 13
rect 177 12 178 13
rect 178 12 179 13
rect 183 12 184 13
rect 184 12 185 13
rect 185 12 186 13
rect 188 12 189 13
rect 189 12 190 13
rect 190 12 191 13
rect 191 12 192 13
rect 196 12 197 13
rect 197 12 198 13
rect 198 12 199 13
rect 199 12 200 13
rect 204 12 205 13
rect 205 12 206 13
rect 206 12 207 13
rect 207 12 208 13
rect 210 12 211 13
rect 211 12 212 13
rect 212 12 213 13
rect 213 12 214 13
rect 221 12 222 13
rect 222 12 223 13
rect 223 12 224 13
rect 224 12 225 13
rect 225 12 226 13
rect 226 12 227 13
rect 227 12 228 13
rect 232 12 233 13
rect 233 12 234 13
rect 234 12 235 13
rect 236 12 237 13
rect 237 12 238 13
rect 238 12 239 13
rect 244 12 245 13
rect 245 12 246 13
rect 246 12 247 13
rect 251 12 252 13
rect 252 12 253 13
rect 253 12 254 13
rect 254 12 255 13
rect 256 12 257 13
rect 257 12 258 13
rect 258 12 259 13
rect 259 12 260 13
rect 260 12 261 13
rect 263 12 264 13
rect 264 12 265 13
rect 267 12 268 13
rect 268 12 269 13
rect 272 12 273 13
rect 273 12 274 13
rect 274 12 275 13
rect 275 12 276 13
rect 276 12 277 13
rect 277 12 278 13
rect 278 12 279 13
rect 279 12 280 13
rect 285 12 286 13
rect 286 12 287 13
rect 287 12 288 13
rect 97 11 98 12
rect 98 11 99 12
rect 99 11 100 12
rect 100 11 101 12
rect 101 11 102 12
rect 102 11 103 12
rect 103 11 104 12
rect 104 11 105 12
rect 123 11 124 12
rect 124 11 125 12
rect 125 11 126 12
rect 126 11 127 12
rect 127 11 128 12
rect 128 11 129 12
rect 129 11 130 12
rect 221 11 222 12
rect 222 11 223 12
rect 223 11 224 12
rect 273 11 274 12
rect 274 11 275 12
rect 275 11 276 12
rect 276 11 277 12
rect 277 11 278 12
rect 278 11 279 12
rect 279 11 280 12
rect 97 10 98 11
rect 98 10 99 11
rect 99 10 100 11
rect 100 10 101 11
rect 101 10 102 11
rect 102 10 103 11
rect 103 10 104 11
rect 104 10 105 11
rect 123 10 124 11
rect 124 10 125 11
rect 125 10 126 11
rect 126 10 127 11
rect 127 10 128 11
rect 128 10 129 11
rect 129 10 130 11
rect 221 10 222 11
rect 222 10 223 11
rect 223 10 224 11
rect 273 10 274 11
rect 274 10 275 11
rect 275 10 276 11
rect 276 10 277 11
rect 277 10 278 11
rect 278 10 279 11
rect 279 10 280 11
rect 97 9 98 10
rect 98 9 99 10
rect 99 9 100 10
rect 100 9 101 10
rect 101 9 102 10
rect 102 9 103 10
rect 103 9 104 10
rect 104 9 105 10
rect 123 9 124 10
rect 124 9 125 10
rect 125 9 126 10
rect 126 9 127 10
rect 127 9 128 10
rect 128 9 129 10
rect 129 9 130 10
rect 221 9 222 10
rect 222 9 223 10
rect 223 9 224 10
rect 273 9 274 10
rect 274 9 275 10
rect 275 9 276 10
rect 276 9 277 10
rect 277 9 278 10
rect 278 9 279 10
rect 279 9 280 10
rect 97 8 98 9
rect 98 8 99 9
rect 99 8 100 9
rect 100 8 101 9
rect 101 8 102 9
rect 102 8 103 9
rect 103 8 104 9
rect 104 8 105 9
rect 123 8 124 9
rect 124 8 125 9
rect 125 8 126 9
rect 126 8 127 9
rect 127 8 128 9
rect 128 8 129 9
rect 129 8 130 9
rect 221 8 222 9
rect 222 8 223 9
rect 223 8 224 9
rect 273 8 274 9
rect 274 8 275 9
rect 275 8 276 9
rect 276 8 277 9
rect 277 8 278 9
rect 278 8 279 9
rect 279 8 280 9
rect 96 7 97 8
rect 97 7 98 8
rect 103 7 104 8
rect 104 7 105 8
rect 122 7 123 8
rect 123 7 124 8
rect 129 7 130 8
rect 221 7 222 8
rect 222 7 223 8
rect 223 7 224 8
rect 272 7 273 8
rect 273 7 274 8
rect 279 7 280 8
rect 96 6 97 7
rect 97 6 98 7
rect 103 6 104 7
rect 104 6 105 7
rect 122 6 123 7
rect 123 6 124 7
rect 129 6 130 7
rect 221 6 222 7
rect 222 6 223 7
rect 223 6 224 7
rect 272 6 273 7
rect 273 6 274 7
rect 279 6 280 7
rect 96 